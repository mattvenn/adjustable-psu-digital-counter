magic
tech sky130A
magscale 1 2
timestamp 1738603755
<< metal2 >>
rect 7264 2753 7444 3324
rect 8912 2783 9092 3244
rect 7260 2583 7269 2753
rect 7439 2583 7448 2753
rect 8908 2613 8917 2783
rect 9087 2613 9096 2783
rect 10594 2753 10774 3258
rect 12226 3209 12406 3310
rect 12222 3039 12231 3209
rect 12401 3039 12410 3209
rect 13858 3143 14038 3346
rect 12226 3034 12406 3039
rect 13854 2973 13863 3143
rect 14033 2973 14042 3143
rect 15540 3091 15720 3318
rect 13858 2968 14038 2973
rect 15536 2921 15545 3091
rect 15715 2921 15724 3091
rect 15540 2916 15720 2921
rect 8912 2608 9092 2613
rect 10590 2583 10599 2753
rect 10769 2583 10778 2753
rect 7264 2578 7444 2583
rect 10594 2578 10774 2583
<< via2 >>
rect 7269 2583 7439 2753
rect 8917 2613 9087 2783
rect 12231 3039 12401 3209
rect 13863 2973 14033 3143
rect 15545 2921 15715 3091
rect 10599 2583 10769 2753
<< metal3 >>
rect 776 16174 1220 16194
rect 776 16173 16936 16174
rect 776 15775 801 16173
rect 1199 15775 16936 16173
rect 776 15774 16936 15775
rect 776 15758 1220 15774
rect 9090 14809 9406 15774
rect 9085 14495 9091 14809
rect 9405 14495 9411 14809
rect 9090 14494 9406 14495
rect 12226 3209 12406 3214
rect 12226 3039 12231 3209
rect 12401 3039 12406 3209
rect 8912 2783 9092 2788
rect 7264 2753 7444 2758
rect 7264 2583 7269 2753
rect 7439 2583 7444 2753
rect 7264 2383 7444 2583
rect 8912 2613 8917 2783
rect 9087 2613 9092 2783
rect 8912 2529 9092 2613
rect 10594 2753 10774 2758
rect 10594 2583 10599 2753
rect 10769 2583 10774 2753
rect 12226 2647 12406 3039
rect 13858 3143 14038 3148
rect 13858 3015 13863 3143
rect 14033 3015 14038 3143
rect 15540 3091 15720 3096
rect 13853 2837 13859 3015
rect 14037 2837 14043 3015
rect 15540 2921 15545 3091
rect 15715 2921 15720 3091
rect 15540 2919 15720 2921
rect 13858 2836 14038 2837
rect 15535 2741 15541 2919
rect 15719 2741 15725 2919
rect 15540 2740 15720 2741
rect 7259 2205 7265 2383
rect 7443 2205 7449 2383
rect 8907 2351 8913 2529
rect 9091 2351 9097 2529
rect 10594 2515 10774 2583
rect 8912 2350 9092 2351
rect 10589 2337 10595 2515
rect 10773 2337 10779 2515
rect 12221 2469 12227 2647
rect 12405 2469 12411 2647
rect 12226 2468 12406 2469
rect 10594 2336 10774 2337
rect 7264 2204 7444 2205
<< via3 >>
rect 801 15775 1199 16173
rect 9091 14495 9405 14809
rect 13859 2973 13863 3015
rect 13863 2973 14033 3015
rect 14033 2973 14037 3015
rect 13859 2837 14037 2973
rect 15541 2741 15719 2919
rect 7265 2205 7443 2383
rect 8913 2351 9091 2529
rect 10595 2337 10773 2515
rect 12227 2469 12405 2647
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 200 1000 600 44152
rect 800 16173 1200 44152
rect 800 15775 801 16173
rect 1199 15775 1200 16173
rect 800 1000 1200 15775
rect 1400 15538 1800 44152
rect 1400 15138 16890 15538
rect 1400 1000 1800 15138
rect 7970 11922 8370 15138
rect 9090 14809 9406 14810
rect 9090 14495 9091 14809
rect 9405 14495 9406 14809
rect 9090 12108 9406 14495
rect 13858 3015 14038 3016
rect 13858 2837 13859 3015
rect 14037 2837 14038 3015
rect 12226 2647 12406 2662
rect 12226 2604 12227 2647
rect 8912 2529 9092 2564
rect 6020 2383 7444 2384
rect 6020 2342 7265 2383
rect 6010 2205 7265 2342
rect 7443 2205 7444 2383
rect 8912 2351 8913 2529
rect 9091 2351 9092 2529
rect 8912 2276 9092 2351
rect 10594 2515 10774 2530
rect 10594 2337 10595 2515
rect 10773 2337 10774 2515
rect 12216 2482 12227 2604
rect 10594 2324 10774 2337
rect 6010 2204 7444 2205
rect 6010 1272 6190 2204
rect 8890 2142 9092 2276
rect 10586 2142 10774 2324
rect 12094 2469 12227 2482
rect 12405 2469 12406 2647
rect 12094 2302 12406 2469
rect 13858 2622 14038 2837
rect 15540 2919 15720 2920
rect 15540 2741 15541 2919
rect 15719 2741 15720 2919
rect 6010 1092 8094 1272
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 1092
rect 8890 334 9070 2142
rect 10586 810 10766 2142
rect 12216 1222 12396 2302
rect 13858 2142 14058 2622
rect 15540 2358 15720 2741
rect 15524 2178 27414 2358
rect 13878 1700 14058 2142
rect 13878 1520 23550 1700
rect 12216 1042 19686 1222
rect 10586 630 15822 810
rect 8890 154 11958 334
rect 11778 0 11958 154
rect 15642 0 15822 630
rect 19506 0 19686 1042
rect 23370 0 23550 1520
rect 27234 0 27414 2178
use count_macro  count_macro_0
timestamp 1738603755
transform 1 0 6486 0 1 3070
box 514 0 9544 9296
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 1600 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
