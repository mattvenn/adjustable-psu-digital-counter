magic
tech sky130A
magscale 1 2
timestamp 1738600851
<< viali >>
rect 4905 2941 4939 2975
rect 5181 2941 5215 2975
rect 6285 2805 6319 2839
rect 3157 2601 3191 2635
rect 4445 2465 4479 2499
rect 7665 2465 7699 2499
rect 8033 2465 8067 2499
rect 5089 2397 5123 2431
rect 7941 2397 7975 2431
rect 8585 2397 8619 2431
rect 5457 2329 5491 2363
rect 5549 2261 5583 2295
rect 6377 2261 6411 2295
rect 4169 1989 4203 2023
rect 2513 1853 2547 1887
rect 3801 1853 3835 1887
rect 3985 1853 4019 1887
rect 4169 1853 4203 1887
rect 8401 1853 8435 1887
rect 8953 1853 8987 1887
rect 6653 1785 6687 1819
rect 3065 1717 3099 1751
rect 3249 1717 3283 1751
rect 5365 1717 5399 1751
rect 7389 1717 7423 1751
rect 2513 1513 2547 1547
rect 5089 1513 5123 1547
rect 6009 1513 6043 1547
rect 7297 1445 7331 1479
rect 8953 1445 8987 1479
rect 2145 1377 2179 1411
rect 2329 1377 2363 1411
rect 3985 1377 4019 1411
rect 4261 1377 4295 1411
rect 5550 1377 5584 1411
rect 6561 1377 6595 1411
rect 6745 1377 6779 1411
rect 7021 1377 7055 1411
rect 8861 1377 8895 1411
rect 2053 1309 2087 1343
rect 4905 1309 4939 1343
rect 5273 1309 5307 1343
rect 5365 1309 5399 1343
rect 5457 1309 5491 1343
rect 5825 1309 5859 1343
rect 5917 1309 5951 1343
rect 6193 1309 6227 1343
rect 6285 1309 6319 1343
rect 6653 1309 6687 1343
rect 2697 1173 2731 1207
rect 4353 1173 4387 1207
rect 6469 1173 6503 1207
rect 8769 1173 8803 1207
rect 2697 969 2731 1003
rect 3065 969 3099 1003
rect 5273 969 5307 1003
rect 5825 969 5859 1003
rect 7941 969 7975 1003
rect 8861 969 8895 1003
rect 3525 833 3559 867
rect 6285 833 6319 867
rect 2421 765 2455 799
rect 2789 765 2823 799
rect 3801 765 3835 799
rect 5457 765 5491 799
rect 6009 765 6043 799
rect 6101 765 6135 799
rect 6193 765 6227 799
rect 6469 765 6503 799
rect 9045 765 9079 799
rect 2697 697 2731 731
rect 3065 697 3099 731
rect 2513 629 2547 663
rect 2881 629 2915 663
rect 4905 629 4939 663
<< metal1 >>
rect 552 9274 9544 9296
rect 552 9222 2606 9274
rect 2658 9222 2670 9274
rect 2722 9222 2734 9274
rect 2786 9222 2798 9274
rect 2850 9222 2862 9274
rect 2914 9222 4814 9274
rect 4866 9222 4878 9274
rect 4930 9222 4942 9274
rect 4994 9222 5006 9274
rect 5058 9222 5070 9274
rect 5122 9222 7022 9274
rect 7074 9222 7086 9274
rect 7138 9222 7150 9274
rect 7202 9222 7214 9274
rect 7266 9222 7278 9274
rect 7330 9222 9230 9274
rect 9282 9222 9294 9274
rect 9346 9222 9358 9274
rect 9410 9222 9422 9274
rect 9474 9222 9486 9274
rect 9538 9222 9544 9274
rect 552 9200 9544 9222
rect 552 8730 9384 8752
rect 552 8678 1502 8730
rect 1554 8678 1566 8730
rect 1618 8678 1630 8730
rect 1682 8678 1694 8730
rect 1746 8678 1758 8730
rect 1810 8678 3710 8730
rect 3762 8678 3774 8730
rect 3826 8678 3838 8730
rect 3890 8678 3902 8730
rect 3954 8678 3966 8730
rect 4018 8678 5918 8730
rect 5970 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 8126 8730
rect 8178 8678 8190 8730
rect 8242 8678 8254 8730
rect 8306 8678 8318 8730
rect 8370 8678 8382 8730
rect 8434 8678 9384 8730
rect 552 8656 9384 8678
rect 552 8186 9544 8208
rect 552 8134 2606 8186
rect 2658 8134 2670 8186
rect 2722 8134 2734 8186
rect 2786 8134 2798 8186
rect 2850 8134 2862 8186
rect 2914 8134 4814 8186
rect 4866 8134 4878 8186
rect 4930 8134 4942 8186
rect 4994 8134 5006 8186
rect 5058 8134 5070 8186
rect 5122 8134 7022 8186
rect 7074 8134 7086 8186
rect 7138 8134 7150 8186
rect 7202 8134 7214 8186
rect 7266 8134 7278 8186
rect 7330 8134 9230 8186
rect 9282 8134 9294 8186
rect 9346 8134 9358 8186
rect 9410 8134 9422 8186
rect 9474 8134 9486 8186
rect 9538 8134 9544 8186
rect 552 8112 9544 8134
rect 552 7642 9384 7664
rect 552 7590 1502 7642
rect 1554 7590 1566 7642
rect 1618 7590 1630 7642
rect 1682 7590 1694 7642
rect 1746 7590 1758 7642
rect 1810 7590 3710 7642
rect 3762 7590 3774 7642
rect 3826 7590 3838 7642
rect 3890 7590 3902 7642
rect 3954 7590 3966 7642
rect 4018 7590 5918 7642
rect 5970 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 8126 7642
rect 8178 7590 8190 7642
rect 8242 7590 8254 7642
rect 8306 7590 8318 7642
rect 8370 7590 8382 7642
rect 8434 7590 9384 7642
rect 552 7568 9384 7590
rect 552 7098 9544 7120
rect 552 7046 2606 7098
rect 2658 7046 2670 7098
rect 2722 7046 2734 7098
rect 2786 7046 2798 7098
rect 2850 7046 2862 7098
rect 2914 7046 4814 7098
rect 4866 7046 4878 7098
rect 4930 7046 4942 7098
rect 4994 7046 5006 7098
rect 5058 7046 5070 7098
rect 5122 7046 7022 7098
rect 7074 7046 7086 7098
rect 7138 7046 7150 7098
rect 7202 7046 7214 7098
rect 7266 7046 7278 7098
rect 7330 7046 9230 7098
rect 9282 7046 9294 7098
rect 9346 7046 9358 7098
rect 9410 7046 9422 7098
rect 9474 7046 9486 7098
rect 9538 7046 9544 7098
rect 552 7024 9544 7046
rect 552 6554 9384 6576
rect 552 6502 1502 6554
rect 1554 6502 1566 6554
rect 1618 6502 1630 6554
rect 1682 6502 1694 6554
rect 1746 6502 1758 6554
rect 1810 6502 3710 6554
rect 3762 6502 3774 6554
rect 3826 6502 3838 6554
rect 3890 6502 3902 6554
rect 3954 6502 3966 6554
rect 4018 6502 5918 6554
rect 5970 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 8126 6554
rect 8178 6502 8190 6554
rect 8242 6502 8254 6554
rect 8306 6502 8318 6554
rect 8370 6502 8382 6554
rect 8434 6502 9384 6554
rect 552 6480 9384 6502
rect 552 6010 9544 6032
rect 552 5958 2606 6010
rect 2658 5958 2670 6010
rect 2722 5958 2734 6010
rect 2786 5958 2798 6010
rect 2850 5958 2862 6010
rect 2914 5958 4814 6010
rect 4866 5958 4878 6010
rect 4930 5958 4942 6010
rect 4994 5958 5006 6010
rect 5058 5958 5070 6010
rect 5122 5958 7022 6010
rect 7074 5958 7086 6010
rect 7138 5958 7150 6010
rect 7202 5958 7214 6010
rect 7266 5958 7278 6010
rect 7330 5958 9230 6010
rect 9282 5958 9294 6010
rect 9346 5958 9358 6010
rect 9410 5958 9422 6010
rect 9474 5958 9486 6010
rect 9538 5958 9544 6010
rect 552 5936 9544 5958
rect 552 5466 9384 5488
rect 552 5414 1502 5466
rect 1554 5414 1566 5466
rect 1618 5414 1630 5466
rect 1682 5414 1694 5466
rect 1746 5414 1758 5466
rect 1810 5414 3710 5466
rect 3762 5414 3774 5466
rect 3826 5414 3838 5466
rect 3890 5414 3902 5466
rect 3954 5414 3966 5466
rect 4018 5414 5918 5466
rect 5970 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 8126 5466
rect 8178 5414 8190 5466
rect 8242 5414 8254 5466
rect 8306 5414 8318 5466
rect 8370 5414 8382 5466
rect 8434 5414 9384 5466
rect 552 5392 9384 5414
rect 552 4922 9544 4944
rect 552 4870 2606 4922
rect 2658 4870 2670 4922
rect 2722 4870 2734 4922
rect 2786 4870 2798 4922
rect 2850 4870 2862 4922
rect 2914 4870 4814 4922
rect 4866 4870 4878 4922
rect 4930 4870 4942 4922
rect 4994 4870 5006 4922
rect 5058 4870 5070 4922
rect 5122 4870 7022 4922
rect 7074 4870 7086 4922
rect 7138 4870 7150 4922
rect 7202 4870 7214 4922
rect 7266 4870 7278 4922
rect 7330 4870 9230 4922
rect 9282 4870 9294 4922
rect 9346 4870 9358 4922
rect 9410 4870 9422 4922
rect 9474 4870 9486 4922
rect 9538 4870 9544 4922
rect 552 4848 9544 4870
rect 552 4378 9384 4400
rect 552 4326 1502 4378
rect 1554 4326 1566 4378
rect 1618 4326 1630 4378
rect 1682 4326 1694 4378
rect 1746 4326 1758 4378
rect 1810 4326 3710 4378
rect 3762 4326 3774 4378
rect 3826 4326 3838 4378
rect 3890 4326 3902 4378
rect 3954 4326 3966 4378
rect 4018 4326 5918 4378
rect 5970 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 8126 4378
rect 8178 4326 8190 4378
rect 8242 4326 8254 4378
rect 8306 4326 8318 4378
rect 8370 4326 8382 4378
rect 8434 4326 9384 4378
rect 552 4304 9384 4326
rect 552 3834 9544 3856
rect 552 3782 2606 3834
rect 2658 3782 2670 3834
rect 2722 3782 2734 3834
rect 2786 3782 2798 3834
rect 2850 3782 2862 3834
rect 2914 3782 4814 3834
rect 4866 3782 4878 3834
rect 4930 3782 4942 3834
rect 4994 3782 5006 3834
rect 5058 3782 5070 3834
rect 5122 3782 7022 3834
rect 7074 3782 7086 3834
rect 7138 3782 7150 3834
rect 7202 3782 7214 3834
rect 7266 3782 7278 3834
rect 7330 3782 9230 3834
rect 9282 3782 9294 3834
rect 9346 3782 9358 3834
rect 9410 3782 9422 3834
rect 9474 3782 9486 3834
rect 9538 3782 9544 3834
rect 552 3760 9544 3782
rect 552 3290 9384 3312
rect 552 3238 1502 3290
rect 1554 3238 1566 3290
rect 1618 3238 1630 3290
rect 1682 3238 1694 3290
rect 1746 3238 1758 3290
rect 1810 3238 3710 3290
rect 3762 3238 3774 3290
rect 3826 3238 3838 3290
rect 3890 3238 3902 3290
rect 3954 3238 3966 3290
rect 4018 3238 5918 3290
rect 5970 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 8126 3290
rect 8178 3238 8190 3290
rect 8242 3238 8254 3290
rect 8306 3238 8318 3290
rect 8370 3238 8382 3290
rect 8434 3238 9384 3290
rect 552 3216 9384 3238
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4212 2944 4905 2972
rect 4212 2932 4218 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 5166 2932 5172 2984
rect 5224 2932 5230 2984
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 6273 2839 6331 2845
rect 6273 2836 6285 2839
rect 5868 2808 6285 2836
rect 5868 2796 5874 2808
rect 6273 2805 6285 2808
rect 6319 2805 6331 2839
rect 6273 2799 6331 2805
rect 552 2746 9544 2768
rect 552 2694 2606 2746
rect 2658 2694 2670 2746
rect 2722 2694 2734 2746
rect 2786 2694 2798 2746
rect 2850 2694 2862 2746
rect 2914 2694 4814 2746
rect 4866 2694 4878 2746
rect 4930 2694 4942 2746
rect 4994 2694 5006 2746
rect 5058 2694 5070 2746
rect 5122 2694 7022 2746
rect 7074 2694 7086 2746
rect 7138 2694 7150 2746
rect 7202 2694 7214 2746
rect 7266 2694 7278 2746
rect 7330 2694 9230 2746
rect 9282 2694 9294 2746
rect 9346 2694 9358 2746
rect 9410 2694 9422 2746
rect 9474 2694 9486 2746
rect 9538 2694 9544 2746
rect 552 2672 9544 2694
rect 3145 2635 3203 2641
rect 3145 2601 3157 2635
rect 3191 2632 3203 2635
rect 4154 2632 4160 2644
rect 3191 2604 4160 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4430 2456 4436 2508
rect 4488 2456 4494 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7699 2468 8033 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8021 2459 8079 2465
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5350 2428 5356 2440
rect 5123 2400 5356 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 5534 2252 5540 2304
rect 5592 2252 5598 2304
rect 6362 2252 6368 2304
rect 6420 2252 6426 2304
rect 552 2202 9384 2224
rect 552 2150 1502 2202
rect 1554 2150 1566 2202
rect 1618 2150 1630 2202
rect 1682 2150 1694 2202
rect 1746 2150 1758 2202
rect 1810 2150 3710 2202
rect 3762 2150 3774 2202
rect 3826 2150 3838 2202
rect 3890 2150 3902 2202
rect 3954 2150 3966 2202
rect 4018 2150 5918 2202
rect 5970 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 8126 2202
rect 8178 2150 8190 2202
rect 8242 2150 8254 2202
rect 8306 2150 8318 2202
rect 8370 2150 8382 2202
rect 8434 2150 9384 2202
rect 552 2128 9384 2150
rect 4157 2023 4215 2029
rect 4157 1989 4169 2023
rect 4203 2020 4215 2023
rect 4246 2020 4252 2032
rect 4203 1992 4252 2020
rect 4203 1989 4215 1992
rect 4157 1983 4215 1989
rect 4246 1980 4252 1992
rect 4304 1980 4310 2032
rect 2498 1844 2504 1896
rect 2556 1844 2562 1896
rect 3786 1844 3792 1896
rect 3844 1844 3850 1896
rect 3973 1887 4031 1893
rect 3973 1853 3985 1887
rect 4019 1853 4031 1887
rect 3973 1847 4031 1853
rect 4157 1887 4215 1893
rect 4157 1853 4169 1887
rect 4203 1884 4215 1887
rect 4706 1884 4712 1896
rect 4203 1856 4712 1884
rect 4203 1853 4215 1856
rect 4157 1847 4215 1853
rect 3418 1776 3424 1828
rect 3476 1816 3482 1828
rect 3988 1816 4016 1847
rect 4706 1844 4712 1856
rect 4764 1844 4770 1896
rect 6730 1844 6736 1896
rect 6788 1884 6794 1896
rect 8389 1887 8447 1893
rect 8389 1884 8401 1887
rect 6788 1856 8401 1884
rect 6788 1844 6794 1856
rect 8389 1853 8401 1856
rect 8435 1853 8447 1887
rect 8389 1847 8447 1853
rect 8938 1844 8944 1896
rect 8996 1844 9002 1896
rect 3476 1788 4016 1816
rect 6641 1819 6699 1825
rect 3476 1776 3482 1788
rect 6641 1785 6653 1819
rect 6687 1816 6699 1819
rect 7466 1816 7472 1828
rect 6687 1788 7472 1816
rect 6687 1785 6699 1788
rect 6641 1779 6699 1785
rect 7466 1776 7472 1788
rect 7524 1776 7530 1828
rect 3050 1708 3056 1760
rect 3108 1708 3114 1760
rect 3234 1708 3240 1760
rect 3292 1708 3298 1760
rect 4430 1708 4436 1760
rect 4488 1748 4494 1760
rect 5353 1751 5411 1757
rect 5353 1748 5365 1751
rect 4488 1720 5365 1748
rect 4488 1708 4494 1720
rect 5353 1717 5365 1720
rect 5399 1748 5411 1751
rect 6454 1748 6460 1760
rect 5399 1720 6460 1748
rect 5399 1717 5411 1720
rect 5353 1711 5411 1717
rect 6454 1708 6460 1720
rect 6512 1708 6518 1760
rect 7374 1708 7380 1760
rect 7432 1708 7438 1760
rect 552 1658 9544 1680
rect 552 1606 2606 1658
rect 2658 1606 2670 1658
rect 2722 1606 2734 1658
rect 2786 1606 2798 1658
rect 2850 1606 2862 1658
rect 2914 1606 4814 1658
rect 4866 1606 4878 1658
rect 4930 1606 4942 1658
rect 4994 1606 5006 1658
rect 5058 1606 5070 1658
rect 5122 1606 7022 1658
rect 7074 1606 7086 1658
rect 7138 1606 7150 1658
rect 7202 1606 7214 1658
rect 7266 1606 7278 1658
rect 7330 1606 9230 1658
rect 9282 1606 9294 1658
rect 9346 1606 9358 1658
rect 9410 1606 9422 1658
rect 9474 1606 9486 1658
rect 9538 1606 9544 1658
rect 552 1584 9544 1606
rect 2498 1504 2504 1556
rect 2556 1504 2562 1556
rect 4706 1504 4712 1556
rect 4764 1544 4770 1556
rect 5077 1547 5135 1553
rect 5077 1544 5089 1547
rect 4764 1516 5089 1544
rect 4764 1504 4770 1516
rect 5077 1513 5089 1516
rect 5123 1513 5135 1547
rect 5997 1547 6055 1553
rect 5997 1544 6009 1547
rect 5077 1507 5135 1513
rect 5276 1516 6009 1544
rect 3234 1476 3240 1488
rect 2148 1448 3240 1476
rect 2148 1417 2176 1448
rect 3234 1436 3240 1448
rect 3292 1436 3298 1488
rect 2133 1411 2191 1417
rect 2133 1377 2145 1411
rect 2179 1377 2191 1411
rect 2133 1371 2191 1377
rect 2314 1368 2320 1420
rect 2372 1368 2378 1420
rect 3050 1368 3056 1420
rect 3108 1408 3114 1420
rect 3973 1411 4031 1417
rect 3973 1408 3985 1411
rect 3108 1380 3985 1408
rect 3108 1368 3114 1380
rect 3973 1377 3985 1380
rect 4019 1377 4031 1411
rect 3973 1371 4031 1377
rect 4154 1368 4160 1420
rect 4212 1408 4218 1420
rect 4249 1411 4307 1417
rect 4249 1408 4261 1411
rect 4212 1380 4261 1408
rect 4212 1368 4218 1380
rect 4249 1377 4261 1380
rect 4295 1377 4307 1411
rect 5276 1408 5304 1516
rect 5997 1513 6009 1516
rect 6043 1544 6055 1547
rect 6270 1544 6276 1556
rect 6043 1516 6276 1544
rect 6043 1513 6055 1516
rect 5997 1507 6055 1513
rect 6270 1504 6276 1516
rect 6328 1504 6334 1556
rect 7926 1544 7932 1556
rect 7024 1516 7932 1544
rect 5538 1411 5596 1417
rect 4249 1371 4307 1377
rect 4816 1380 5396 1408
rect 1302 1300 1308 1352
rect 1360 1340 1366 1352
rect 2041 1343 2099 1349
rect 2041 1340 2053 1343
rect 1360 1312 2053 1340
rect 1360 1300 1366 1312
rect 2041 1309 2053 1312
rect 2087 1309 2099 1343
rect 2041 1303 2099 1309
rect 4816 1272 4844 1380
rect 4890 1300 4896 1352
rect 4948 1340 4954 1352
rect 5368 1349 5396 1380
rect 5538 1377 5550 1411
rect 5584 1408 5596 1411
rect 5626 1408 5632 1420
rect 5584 1380 5632 1408
rect 5584 1377 5596 1380
rect 5538 1371 5596 1377
rect 5626 1368 5632 1380
rect 5684 1368 5690 1420
rect 6362 1408 6368 1420
rect 5736 1380 6368 1408
rect 5736 1352 5764 1380
rect 5261 1343 5319 1349
rect 5261 1340 5273 1343
rect 4948 1312 5273 1340
rect 4948 1300 4954 1312
rect 5261 1309 5273 1312
rect 5307 1309 5319 1343
rect 5261 1303 5319 1309
rect 5353 1343 5411 1349
rect 5353 1309 5365 1343
rect 5399 1309 5411 1343
rect 5353 1303 5411 1309
rect 5445 1343 5503 1349
rect 5445 1309 5457 1343
rect 5491 1340 5503 1343
rect 5718 1340 5724 1352
rect 5491 1312 5724 1340
rect 5491 1309 5503 1312
rect 5445 1303 5503 1309
rect 4264 1244 4844 1272
rect 5276 1272 5304 1303
rect 5718 1300 5724 1312
rect 5776 1300 5782 1352
rect 5810 1300 5816 1352
rect 5868 1300 5874 1352
rect 6196 1349 6224 1380
rect 6362 1368 6368 1380
rect 6420 1408 6426 1420
rect 6549 1411 6607 1417
rect 6549 1408 6561 1411
rect 6420 1380 6561 1408
rect 6420 1368 6426 1380
rect 6549 1377 6561 1380
rect 6595 1377 6607 1411
rect 6549 1371 6607 1377
rect 6730 1368 6736 1420
rect 6788 1368 6794 1420
rect 7024 1417 7052 1516
rect 7926 1504 7932 1516
rect 7984 1504 7990 1556
rect 7285 1479 7343 1485
rect 7285 1445 7297 1479
rect 7331 1476 7343 1479
rect 7374 1476 7380 1488
rect 7331 1448 7380 1476
rect 7331 1445 7343 1448
rect 7285 1439 7343 1445
rect 7374 1436 7380 1448
rect 7432 1436 7438 1488
rect 8941 1479 8999 1485
rect 8941 1476 8953 1479
rect 8510 1448 8953 1476
rect 8941 1445 8953 1448
rect 8987 1445 8999 1479
rect 8941 1439 8999 1445
rect 7009 1411 7067 1417
rect 7009 1377 7021 1411
rect 7055 1377 7067 1411
rect 7009 1371 7067 1377
rect 8846 1368 8852 1420
rect 8904 1368 8910 1420
rect 5905 1343 5963 1349
rect 5905 1309 5917 1343
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6181 1343 6239 1349
rect 6181 1309 6193 1343
rect 6227 1309 6239 1343
rect 6181 1303 6239 1309
rect 6273 1343 6331 1349
rect 6273 1309 6285 1343
rect 6319 1309 6331 1343
rect 6273 1303 6331 1309
rect 6641 1343 6699 1349
rect 6641 1309 6653 1343
rect 6687 1340 6699 1343
rect 8570 1340 8576 1352
rect 6687 1312 8576 1340
rect 6687 1309 6699 1312
rect 6641 1303 6699 1309
rect 5920 1272 5948 1303
rect 5276 1244 5948 1272
rect 6288 1272 6316 1303
rect 8570 1300 8576 1312
rect 8628 1300 8634 1352
rect 6288 1244 6914 1272
rect 2498 1164 2504 1216
rect 2556 1204 2562 1216
rect 2685 1207 2743 1213
rect 2685 1204 2697 1207
rect 2556 1176 2697 1204
rect 2556 1164 2562 1176
rect 2685 1173 2697 1176
rect 2731 1204 2743 1207
rect 3786 1204 3792 1216
rect 2731 1176 3792 1204
rect 2731 1173 2743 1176
rect 2685 1167 2743 1173
rect 3786 1164 3792 1176
rect 3844 1204 3850 1216
rect 4264 1204 4292 1244
rect 3844 1176 4292 1204
rect 4341 1207 4399 1213
rect 3844 1164 3850 1176
rect 4341 1173 4353 1207
rect 4387 1204 4399 1207
rect 4430 1204 4436 1216
rect 4387 1176 4436 1204
rect 4387 1173 4399 1176
rect 4341 1167 4399 1173
rect 4430 1164 4436 1176
rect 4488 1164 4494 1216
rect 5350 1164 5356 1216
rect 5408 1204 5414 1216
rect 6457 1207 6515 1213
rect 6457 1204 6469 1207
rect 5408 1176 6469 1204
rect 5408 1164 5414 1176
rect 6457 1173 6469 1176
rect 6503 1173 6515 1207
rect 6886 1204 6914 1244
rect 8757 1207 8815 1213
rect 8757 1204 8769 1207
rect 6886 1176 8769 1204
rect 6457 1167 6515 1173
rect 8757 1173 8769 1176
rect 8803 1204 8815 1207
rect 8938 1204 8944 1216
rect 8803 1176 8944 1204
rect 8803 1173 8815 1176
rect 8757 1167 8815 1173
rect 8938 1164 8944 1176
rect 8996 1164 9002 1216
rect 552 1114 9384 1136
rect 552 1062 1502 1114
rect 1554 1062 1566 1114
rect 1618 1062 1630 1114
rect 1682 1062 1694 1114
rect 1746 1062 1758 1114
rect 1810 1062 3710 1114
rect 3762 1062 3774 1114
rect 3826 1062 3838 1114
rect 3890 1062 3902 1114
rect 3954 1062 3966 1114
rect 4018 1062 5918 1114
rect 5970 1062 5982 1114
rect 6034 1062 6046 1114
rect 6098 1062 6110 1114
rect 6162 1062 6174 1114
rect 6226 1062 8126 1114
rect 8178 1062 8190 1114
rect 8242 1062 8254 1114
rect 8306 1062 8318 1114
rect 8370 1062 8382 1114
rect 8434 1062 9384 1114
rect 552 1040 9384 1062
rect 2314 960 2320 1012
rect 2372 1000 2378 1012
rect 2685 1003 2743 1009
rect 2685 1000 2697 1003
rect 2372 972 2697 1000
rect 2372 960 2378 972
rect 2685 969 2697 972
rect 2731 969 2743 1003
rect 2685 963 2743 969
rect 3053 1003 3111 1009
rect 3053 969 3065 1003
rect 3099 1000 3111 1003
rect 3418 1000 3424 1012
rect 3099 972 3424 1000
rect 3099 969 3111 972
rect 3053 963 3111 969
rect 3418 960 3424 972
rect 3476 960 3482 1012
rect 3528 972 5120 1000
rect 3528 932 3556 972
rect 2976 904 3556 932
rect 5092 932 5120 972
rect 5166 960 5172 1012
rect 5224 1000 5230 1012
rect 5261 1003 5319 1009
rect 5261 1000 5273 1003
rect 5224 972 5273 1000
rect 5224 960 5230 972
rect 5261 969 5273 972
rect 5307 969 5319 1003
rect 5261 963 5319 969
rect 5442 960 5448 1012
rect 5500 1000 5506 1012
rect 5813 1003 5871 1009
rect 5813 1000 5825 1003
rect 5500 972 5825 1000
rect 5500 960 5506 972
rect 5813 969 5825 972
rect 5859 969 5871 1003
rect 5813 963 5871 969
rect 7926 960 7932 1012
rect 7984 960 7990 1012
rect 8846 960 8852 1012
rect 8904 960 8910 1012
rect 5626 932 5632 944
rect 5092 904 5632 932
rect 2409 799 2467 805
rect 2409 765 2421 799
rect 2455 796 2467 799
rect 2498 796 2504 808
rect 2455 768 2504 796
rect 2455 765 2467 768
rect 2409 759 2467 765
rect 2498 756 2504 768
rect 2556 796 2562 808
rect 2777 799 2835 805
rect 2777 796 2789 799
rect 2556 768 2789 796
rect 2556 756 2562 768
rect 2777 765 2789 768
rect 2823 765 2835 799
rect 2777 759 2835 765
rect 2685 731 2743 737
rect 2685 697 2697 731
rect 2731 728 2743 731
rect 2976 728 3004 904
rect 5626 892 5632 904
rect 5684 932 5690 944
rect 6730 932 6736 944
rect 5684 904 6736 932
rect 5684 892 5690 904
rect 6730 892 6736 904
rect 6788 892 6794 944
rect 3513 867 3571 873
rect 3513 833 3525 867
rect 3559 864 3571 867
rect 4154 864 4160 876
rect 3559 836 4160 864
rect 3559 833 3571 836
rect 3513 827 3571 833
rect 4154 824 4160 836
rect 4212 824 4218 876
rect 5810 824 5816 876
rect 5868 864 5874 876
rect 6273 867 6331 873
rect 6273 864 6285 867
rect 5868 836 6285 864
rect 5868 824 5874 836
rect 6273 833 6285 836
rect 6319 833 6331 867
rect 6273 827 6331 833
rect 3789 799 3847 805
rect 3789 765 3801 799
rect 3835 796 3847 799
rect 4246 796 4252 808
rect 3835 768 4252 796
rect 3835 765 3847 768
rect 3789 759 3847 765
rect 4246 756 4252 768
rect 4304 756 4310 808
rect 5445 799 5503 805
rect 5445 765 5457 799
rect 5491 796 5503 799
rect 5534 796 5540 808
rect 5491 768 5540 796
rect 5491 765 5503 768
rect 5445 759 5503 765
rect 5534 756 5540 768
rect 5592 756 5598 808
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 6089 799 6147 805
rect 6089 765 6101 799
rect 6135 765 6147 799
rect 6089 759 6147 765
rect 6181 799 6239 805
rect 6181 765 6193 799
rect 6227 796 6239 799
rect 6362 796 6368 808
rect 6227 768 6368 796
rect 6227 765 6239 768
rect 6181 759 6239 765
rect 2731 700 3004 728
rect 3053 731 3111 737
rect 2731 697 2743 700
rect 2685 691 2743 697
rect 3053 697 3065 731
rect 3099 697 3111 731
rect 6012 728 6040 759
rect 3053 691 3111 697
rect 4908 700 6040 728
rect 6104 728 6132 759
rect 6362 756 6368 768
rect 6420 756 6426 808
rect 6454 756 6460 808
rect 6512 756 6518 808
rect 9033 799 9091 805
rect 9033 765 9045 799
rect 9079 796 9091 799
rect 9122 796 9128 808
rect 9079 768 9128 796
rect 9079 765 9091 768
rect 9033 759 9091 765
rect 9122 756 9128 768
rect 9180 756 9186 808
rect 6270 728 6276 740
rect 6104 700 6276 728
rect 842 620 848 672
rect 900 660 906 672
rect 1302 660 1308 672
rect 900 632 1308 660
rect 900 620 906 632
rect 1302 620 1308 632
rect 1360 660 1366 672
rect 2501 663 2559 669
rect 2501 660 2513 663
rect 1360 632 2513 660
rect 1360 620 1366 632
rect 2501 629 2513 632
rect 2547 660 2559 663
rect 2869 663 2927 669
rect 2869 660 2881 663
rect 2547 632 2881 660
rect 2547 629 2559 632
rect 2501 623 2559 629
rect 2869 629 2881 632
rect 2915 660 2927 663
rect 2958 660 2964 672
rect 2915 632 2964 660
rect 2915 629 2927 632
rect 2869 623 2927 629
rect 2958 620 2964 632
rect 3016 620 3022 672
rect 3068 660 3096 691
rect 4908 672 4936 700
rect 6270 688 6276 700
rect 6328 688 6334 740
rect 4430 660 4436 672
rect 3068 632 4436 660
rect 4430 620 4436 632
rect 4488 620 4494 672
rect 4522 620 4528 672
rect 4580 660 4586 672
rect 4890 660 4896 672
rect 4580 632 4896 660
rect 4580 620 4586 632
rect 4890 620 4896 632
rect 4948 620 4954 672
rect 552 570 9544 592
rect 552 518 2606 570
rect 2658 518 2670 570
rect 2722 518 2734 570
rect 2786 518 2798 570
rect 2850 518 2862 570
rect 2914 518 4814 570
rect 4866 518 4878 570
rect 4930 518 4942 570
rect 4994 518 5006 570
rect 5058 518 5070 570
rect 5122 518 7022 570
rect 7074 518 7086 570
rect 7138 518 7150 570
rect 7202 518 7214 570
rect 7266 518 7278 570
rect 7330 518 9230 570
rect 9282 518 9294 570
rect 9346 518 9358 570
rect 9410 518 9422 570
rect 9474 518 9486 570
rect 9538 518 9544 570
rect 552 496 9544 518
rect 2958 416 2964 468
rect 3016 456 3022 468
rect 5718 456 5724 468
rect 3016 428 5724 456
rect 3016 416 3022 428
rect 5718 416 5724 428
rect 5776 416 5782 468
<< via1 >>
rect 2606 9222 2658 9274
rect 2670 9222 2722 9274
rect 2734 9222 2786 9274
rect 2798 9222 2850 9274
rect 2862 9222 2914 9274
rect 4814 9222 4866 9274
rect 4878 9222 4930 9274
rect 4942 9222 4994 9274
rect 5006 9222 5058 9274
rect 5070 9222 5122 9274
rect 7022 9222 7074 9274
rect 7086 9222 7138 9274
rect 7150 9222 7202 9274
rect 7214 9222 7266 9274
rect 7278 9222 7330 9274
rect 9230 9222 9282 9274
rect 9294 9222 9346 9274
rect 9358 9222 9410 9274
rect 9422 9222 9474 9274
rect 9486 9222 9538 9274
rect 1502 8678 1554 8730
rect 1566 8678 1618 8730
rect 1630 8678 1682 8730
rect 1694 8678 1746 8730
rect 1758 8678 1810 8730
rect 3710 8678 3762 8730
rect 3774 8678 3826 8730
rect 3838 8678 3890 8730
rect 3902 8678 3954 8730
rect 3966 8678 4018 8730
rect 5918 8678 5970 8730
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 8126 8678 8178 8730
rect 8190 8678 8242 8730
rect 8254 8678 8306 8730
rect 8318 8678 8370 8730
rect 8382 8678 8434 8730
rect 2606 8134 2658 8186
rect 2670 8134 2722 8186
rect 2734 8134 2786 8186
rect 2798 8134 2850 8186
rect 2862 8134 2914 8186
rect 4814 8134 4866 8186
rect 4878 8134 4930 8186
rect 4942 8134 4994 8186
rect 5006 8134 5058 8186
rect 5070 8134 5122 8186
rect 7022 8134 7074 8186
rect 7086 8134 7138 8186
rect 7150 8134 7202 8186
rect 7214 8134 7266 8186
rect 7278 8134 7330 8186
rect 9230 8134 9282 8186
rect 9294 8134 9346 8186
rect 9358 8134 9410 8186
rect 9422 8134 9474 8186
rect 9486 8134 9538 8186
rect 1502 7590 1554 7642
rect 1566 7590 1618 7642
rect 1630 7590 1682 7642
rect 1694 7590 1746 7642
rect 1758 7590 1810 7642
rect 3710 7590 3762 7642
rect 3774 7590 3826 7642
rect 3838 7590 3890 7642
rect 3902 7590 3954 7642
rect 3966 7590 4018 7642
rect 5918 7590 5970 7642
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 8126 7590 8178 7642
rect 8190 7590 8242 7642
rect 8254 7590 8306 7642
rect 8318 7590 8370 7642
rect 8382 7590 8434 7642
rect 2606 7046 2658 7098
rect 2670 7046 2722 7098
rect 2734 7046 2786 7098
rect 2798 7046 2850 7098
rect 2862 7046 2914 7098
rect 4814 7046 4866 7098
rect 4878 7046 4930 7098
rect 4942 7046 4994 7098
rect 5006 7046 5058 7098
rect 5070 7046 5122 7098
rect 7022 7046 7074 7098
rect 7086 7046 7138 7098
rect 7150 7046 7202 7098
rect 7214 7046 7266 7098
rect 7278 7046 7330 7098
rect 9230 7046 9282 7098
rect 9294 7046 9346 7098
rect 9358 7046 9410 7098
rect 9422 7046 9474 7098
rect 9486 7046 9538 7098
rect 1502 6502 1554 6554
rect 1566 6502 1618 6554
rect 1630 6502 1682 6554
rect 1694 6502 1746 6554
rect 1758 6502 1810 6554
rect 3710 6502 3762 6554
rect 3774 6502 3826 6554
rect 3838 6502 3890 6554
rect 3902 6502 3954 6554
rect 3966 6502 4018 6554
rect 5918 6502 5970 6554
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 8126 6502 8178 6554
rect 8190 6502 8242 6554
rect 8254 6502 8306 6554
rect 8318 6502 8370 6554
rect 8382 6502 8434 6554
rect 2606 5958 2658 6010
rect 2670 5958 2722 6010
rect 2734 5958 2786 6010
rect 2798 5958 2850 6010
rect 2862 5958 2914 6010
rect 4814 5958 4866 6010
rect 4878 5958 4930 6010
rect 4942 5958 4994 6010
rect 5006 5958 5058 6010
rect 5070 5958 5122 6010
rect 7022 5958 7074 6010
rect 7086 5958 7138 6010
rect 7150 5958 7202 6010
rect 7214 5958 7266 6010
rect 7278 5958 7330 6010
rect 9230 5958 9282 6010
rect 9294 5958 9346 6010
rect 9358 5958 9410 6010
rect 9422 5958 9474 6010
rect 9486 5958 9538 6010
rect 1502 5414 1554 5466
rect 1566 5414 1618 5466
rect 1630 5414 1682 5466
rect 1694 5414 1746 5466
rect 1758 5414 1810 5466
rect 3710 5414 3762 5466
rect 3774 5414 3826 5466
rect 3838 5414 3890 5466
rect 3902 5414 3954 5466
rect 3966 5414 4018 5466
rect 5918 5414 5970 5466
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 8126 5414 8178 5466
rect 8190 5414 8242 5466
rect 8254 5414 8306 5466
rect 8318 5414 8370 5466
rect 8382 5414 8434 5466
rect 2606 4870 2658 4922
rect 2670 4870 2722 4922
rect 2734 4870 2786 4922
rect 2798 4870 2850 4922
rect 2862 4870 2914 4922
rect 4814 4870 4866 4922
rect 4878 4870 4930 4922
rect 4942 4870 4994 4922
rect 5006 4870 5058 4922
rect 5070 4870 5122 4922
rect 7022 4870 7074 4922
rect 7086 4870 7138 4922
rect 7150 4870 7202 4922
rect 7214 4870 7266 4922
rect 7278 4870 7330 4922
rect 9230 4870 9282 4922
rect 9294 4870 9346 4922
rect 9358 4870 9410 4922
rect 9422 4870 9474 4922
rect 9486 4870 9538 4922
rect 1502 4326 1554 4378
rect 1566 4326 1618 4378
rect 1630 4326 1682 4378
rect 1694 4326 1746 4378
rect 1758 4326 1810 4378
rect 3710 4326 3762 4378
rect 3774 4326 3826 4378
rect 3838 4326 3890 4378
rect 3902 4326 3954 4378
rect 3966 4326 4018 4378
rect 5918 4326 5970 4378
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 8126 4326 8178 4378
rect 8190 4326 8242 4378
rect 8254 4326 8306 4378
rect 8318 4326 8370 4378
rect 8382 4326 8434 4378
rect 2606 3782 2658 3834
rect 2670 3782 2722 3834
rect 2734 3782 2786 3834
rect 2798 3782 2850 3834
rect 2862 3782 2914 3834
rect 4814 3782 4866 3834
rect 4878 3782 4930 3834
rect 4942 3782 4994 3834
rect 5006 3782 5058 3834
rect 5070 3782 5122 3834
rect 7022 3782 7074 3834
rect 7086 3782 7138 3834
rect 7150 3782 7202 3834
rect 7214 3782 7266 3834
rect 7278 3782 7330 3834
rect 9230 3782 9282 3834
rect 9294 3782 9346 3834
rect 9358 3782 9410 3834
rect 9422 3782 9474 3834
rect 9486 3782 9538 3834
rect 1502 3238 1554 3290
rect 1566 3238 1618 3290
rect 1630 3238 1682 3290
rect 1694 3238 1746 3290
rect 1758 3238 1810 3290
rect 3710 3238 3762 3290
rect 3774 3238 3826 3290
rect 3838 3238 3890 3290
rect 3902 3238 3954 3290
rect 3966 3238 4018 3290
rect 5918 3238 5970 3290
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 8126 3238 8178 3290
rect 8190 3238 8242 3290
rect 8254 3238 8306 3290
rect 8318 3238 8370 3290
rect 8382 3238 8434 3290
rect 4160 2932 4212 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 5816 2796 5868 2848
rect 2606 2694 2658 2746
rect 2670 2694 2722 2746
rect 2734 2694 2786 2746
rect 2798 2694 2850 2746
rect 2862 2694 2914 2746
rect 4814 2694 4866 2746
rect 4878 2694 4930 2746
rect 4942 2694 4994 2746
rect 5006 2694 5058 2746
rect 5070 2694 5122 2746
rect 7022 2694 7074 2746
rect 7086 2694 7138 2746
rect 7150 2694 7202 2746
rect 7214 2694 7266 2746
rect 7278 2694 7330 2746
rect 9230 2694 9282 2746
rect 9294 2694 9346 2746
rect 9358 2694 9410 2746
rect 9422 2694 9474 2746
rect 9486 2694 9538 2746
rect 4160 2592 4212 2644
rect 4436 2499 4488 2508
rect 4436 2465 4445 2499
rect 4445 2465 4479 2499
rect 4479 2465 4488 2499
rect 4436 2456 4488 2465
rect 5356 2388 5408 2440
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 5540 2295 5592 2304
rect 5540 2261 5549 2295
rect 5549 2261 5583 2295
rect 5583 2261 5592 2295
rect 5540 2252 5592 2261
rect 6368 2295 6420 2304
rect 6368 2261 6377 2295
rect 6377 2261 6411 2295
rect 6411 2261 6420 2295
rect 6368 2252 6420 2261
rect 1502 2150 1554 2202
rect 1566 2150 1618 2202
rect 1630 2150 1682 2202
rect 1694 2150 1746 2202
rect 1758 2150 1810 2202
rect 3710 2150 3762 2202
rect 3774 2150 3826 2202
rect 3838 2150 3890 2202
rect 3902 2150 3954 2202
rect 3966 2150 4018 2202
rect 5918 2150 5970 2202
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 8126 2150 8178 2202
rect 8190 2150 8242 2202
rect 8254 2150 8306 2202
rect 8318 2150 8370 2202
rect 8382 2150 8434 2202
rect 4252 1980 4304 2032
rect 2504 1887 2556 1896
rect 2504 1853 2513 1887
rect 2513 1853 2547 1887
rect 2547 1853 2556 1887
rect 2504 1844 2556 1853
rect 3792 1887 3844 1896
rect 3792 1853 3801 1887
rect 3801 1853 3835 1887
rect 3835 1853 3844 1887
rect 3792 1844 3844 1853
rect 3424 1776 3476 1828
rect 4712 1844 4764 1896
rect 6736 1844 6788 1896
rect 8944 1887 8996 1896
rect 8944 1853 8953 1887
rect 8953 1853 8987 1887
rect 8987 1853 8996 1887
rect 8944 1844 8996 1853
rect 7472 1776 7524 1828
rect 3056 1751 3108 1760
rect 3056 1717 3065 1751
rect 3065 1717 3099 1751
rect 3099 1717 3108 1751
rect 3056 1708 3108 1717
rect 3240 1751 3292 1760
rect 3240 1717 3249 1751
rect 3249 1717 3283 1751
rect 3283 1717 3292 1751
rect 3240 1708 3292 1717
rect 4436 1708 4488 1760
rect 6460 1708 6512 1760
rect 7380 1751 7432 1760
rect 7380 1717 7389 1751
rect 7389 1717 7423 1751
rect 7423 1717 7432 1751
rect 7380 1708 7432 1717
rect 2606 1606 2658 1658
rect 2670 1606 2722 1658
rect 2734 1606 2786 1658
rect 2798 1606 2850 1658
rect 2862 1606 2914 1658
rect 4814 1606 4866 1658
rect 4878 1606 4930 1658
rect 4942 1606 4994 1658
rect 5006 1606 5058 1658
rect 5070 1606 5122 1658
rect 7022 1606 7074 1658
rect 7086 1606 7138 1658
rect 7150 1606 7202 1658
rect 7214 1606 7266 1658
rect 7278 1606 7330 1658
rect 9230 1606 9282 1658
rect 9294 1606 9346 1658
rect 9358 1606 9410 1658
rect 9422 1606 9474 1658
rect 9486 1606 9538 1658
rect 2504 1547 2556 1556
rect 2504 1513 2513 1547
rect 2513 1513 2547 1547
rect 2547 1513 2556 1547
rect 2504 1504 2556 1513
rect 4712 1504 4764 1556
rect 3240 1436 3292 1488
rect 2320 1411 2372 1420
rect 2320 1377 2329 1411
rect 2329 1377 2363 1411
rect 2363 1377 2372 1411
rect 2320 1368 2372 1377
rect 3056 1368 3108 1420
rect 4160 1368 4212 1420
rect 6276 1504 6328 1556
rect 1308 1300 1360 1352
rect 4896 1343 4948 1352
rect 4896 1309 4905 1343
rect 4905 1309 4939 1343
rect 4939 1309 4948 1343
rect 5632 1368 5684 1420
rect 4896 1300 4948 1309
rect 5724 1300 5776 1352
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 6368 1368 6420 1420
rect 6736 1411 6788 1420
rect 6736 1377 6745 1411
rect 6745 1377 6779 1411
rect 6779 1377 6788 1411
rect 6736 1368 6788 1377
rect 7932 1504 7984 1556
rect 7380 1436 7432 1488
rect 8852 1411 8904 1420
rect 8852 1377 8861 1411
rect 8861 1377 8895 1411
rect 8895 1377 8904 1411
rect 8852 1368 8904 1377
rect 8576 1300 8628 1352
rect 2504 1164 2556 1216
rect 3792 1164 3844 1216
rect 4436 1164 4488 1216
rect 5356 1164 5408 1216
rect 8944 1164 8996 1216
rect 1502 1062 1554 1114
rect 1566 1062 1618 1114
rect 1630 1062 1682 1114
rect 1694 1062 1746 1114
rect 1758 1062 1810 1114
rect 3710 1062 3762 1114
rect 3774 1062 3826 1114
rect 3838 1062 3890 1114
rect 3902 1062 3954 1114
rect 3966 1062 4018 1114
rect 5918 1062 5970 1114
rect 5982 1062 6034 1114
rect 6046 1062 6098 1114
rect 6110 1062 6162 1114
rect 6174 1062 6226 1114
rect 8126 1062 8178 1114
rect 8190 1062 8242 1114
rect 8254 1062 8306 1114
rect 8318 1062 8370 1114
rect 8382 1062 8434 1114
rect 2320 960 2372 1012
rect 3424 960 3476 1012
rect 5172 960 5224 1012
rect 5448 960 5500 1012
rect 7932 1003 7984 1012
rect 7932 969 7941 1003
rect 7941 969 7975 1003
rect 7975 969 7984 1003
rect 7932 960 7984 969
rect 8852 1003 8904 1012
rect 8852 969 8861 1003
rect 8861 969 8895 1003
rect 8895 969 8904 1003
rect 8852 960 8904 969
rect 2504 756 2556 808
rect 5632 892 5684 944
rect 6736 892 6788 944
rect 4160 824 4212 876
rect 5816 824 5868 876
rect 4252 756 4304 808
rect 5540 756 5592 808
rect 6368 756 6420 808
rect 6460 799 6512 808
rect 6460 765 6469 799
rect 6469 765 6503 799
rect 6503 765 6512 799
rect 6460 756 6512 765
rect 9128 756 9180 808
rect 848 620 900 672
rect 1308 620 1360 672
rect 2964 620 3016 672
rect 6276 688 6328 740
rect 4436 620 4488 672
rect 4528 620 4580 672
rect 4896 663 4948 672
rect 4896 629 4905 663
rect 4905 629 4939 663
rect 4939 629 4948 663
rect 4896 620 4948 629
rect 2606 518 2658 570
rect 2670 518 2722 570
rect 2734 518 2786 570
rect 2798 518 2850 570
rect 2862 518 2914 570
rect 4814 518 4866 570
rect 4878 518 4930 570
rect 4942 518 4994 570
rect 5006 518 5058 570
rect 5070 518 5122 570
rect 7022 518 7074 570
rect 7086 518 7138 570
rect 7150 518 7202 570
rect 7214 518 7266 570
rect 7278 518 7330 570
rect 9230 518 9282 570
rect 9294 518 9346 570
rect 9358 518 9410 570
rect 9422 518 9474 570
rect 9486 518 9538 570
rect 2964 416 3016 468
rect 5724 416 5776 468
<< metal2 >>
rect 2606 9276 2914 9285
rect 2606 9274 2612 9276
rect 2668 9274 2692 9276
rect 2748 9274 2772 9276
rect 2828 9274 2852 9276
rect 2908 9274 2914 9276
rect 2668 9222 2670 9274
rect 2850 9222 2852 9274
rect 2606 9220 2612 9222
rect 2668 9220 2692 9222
rect 2748 9220 2772 9222
rect 2828 9220 2852 9222
rect 2908 9220 2914 9222
rect 2606 9211 2914 9220
rect 4814 9276 5122 9285
rect 4814 9274 4820 9276
rect 4876 9274 4900 9276
rect 4956 9274 4980 9276
rect 5036 9274 5060 9276
rect 5116 9274 5122 9276
rect 4876 9222 4878 9274
rect 5058 9222 5060 9274
rect 4814 9220 4820 9222
rect 4876 9220 4900 9222
rect 4956 9220 4980 9222
rect 5036 9220 5060 9222
rect 5116 9220 5122 9222
rect 4814 9211 5122 9220
rect 7022 9276 7330 9285
rect 7022 9274 7028 9276
rect 7084 9274 7108 9276
rect 7164 9274 7188 9276
rect 7244 9274 7268 9276
rect 7324 9274 7330 9276
rect 7084 9222 7086 9274
rect 7266 9222 7268 9274
rect 7022 9220 7028 9222
rect 7084 9220 7108 9222
rect 7164 9220 7188 9222
rect 7244 9220 7268 9222
rect 7324 9220 7330 9222
rect 7022 9211 7330 9220
rect 9230 9276 9538 9285
rect 9230 9274 9236 9276
rect 9292 9274 9316 9276
rect 9372 9274 9396 9276
rect 9452 9274 9476 9276
rect 9532 9274 9538 9276
rect 9292 9222 9294 9274
rect 9474 9222 9476 9274
rect 9230 9220 9236 9222
rect 9292 9220 9316 9222
rect 9372 9220 9396 9222
rect 9452 9220 9476 9222
rect 9532 9220 9538 9222
rect 9230 9211 9538 9220
rect 1502 8732 1810 8741
rect 1502 8730 1508 8732
rect 1564 8730 1588 8732
rect 1644 8730 1668 8732
rect 1724 8730 1748 8732
rect 1804 8730 1810 8732
rect 1564 8678 1566 8730
rect 1746 8678 1748 8730
rect 1502 8676 1508 8678
rect 1564 8676 1588 8678
rect 1644 8676 1668 8678
rect 1724 8676 1748 8678
rect 1804 8676 1810 8678
rect 1502 8667 1810 8676
rect 3710 8732 4018 8741
rect 3710 8730 3716 8732
rect 3772 8730 3796 8732
rect 3852 8730 3876 8732
rect 3932 8730 3956 8732
rect 4012 8730 4018 8732
rect 3772 8678 3774 8730
rect 3954 8678 3956 8730
rect 3710 8676 3716 8678
rect 3772 8676 3796 8678
rect 3852 8676 3876 8678
rect 3932 8676 3956 8678
rect 4012 8676 4018 8678
rect 3710 8667 4018 8676
rect 5918 8732 6226 8741
rect 5918 8730 5924 8732
rect 5980 8730 6004 8732
rect 6060 8730 6084 8732
rect 6140 8730 6164 8732
rect 6220 8730 6226 8732
rect 5980 8678 5982 8730
rect 6162 8678 6164 8730
rect 5918 8676 5924 8678
rect 5980 8676 6004 8678
rect 6060 8676 6084 8678
rect 6140 8676 6164 8678
rect 6220 8676 6226 8678
rect 5918 8667 6226 8676
rect 8126 8732 8434 8741
rect 8126 8730 8132 8732
rect 8188 8730 8212 8732
rect 8268 8730 8292 8732
rect 8348 8730 8372 8732
rect 8428 8730 8434 8732
rect 8188 8678 8190 8730
rect 8370 8678 8372 8730
rect 8126 8676 8132 8678
rect 8188 8676 8212 8678
rect 8268 8676 8292 8678
rect 8348 8676 8372 8678
rect 8428 8676 8434 8678
rect 8126 8667 8434 8676
rect 2606 8188 2914 8197
rect 2606 8186 2612 8188
rect 2668 8186 2692 8188
rect 2748 8186 2772 8188
rect 2828 8186 2852 8188
rect 2908 8186 2914 8188
rect 2668 8134 2670 8186
rect 2850 8134 2852 8186
rect 2606 8132 2612 8134
rect 2668 8132 2692 8134
rect 2748 8132 2772 8134
rect 2828 8132 2852 8134
rect 2908 8132 2914 8134
rect 2606 8123 2914 8132
rect 4814 8188 5122 8197
rect 4814 8186 4820 8188
rect 4876 8186 4900 8188
rect 4956 8186 4980 8188
rect 5036 8186 5060 8188
rect 5116 8186 5122 8188
rect 4876 8134 4878 8186
rect 5058 8134 5060 8186
rect 4814 8132 4820 8134
rect 4876 8132 4900 8134
rect 4956 8132 4980 8134
rect 5036 8132 5060 8134
rect 5116 8132 5122 8134
rect 4814 8123 5122 8132
rect 7022 8188 7330 8197
rect 7022 8186 7028 8188
rect 7084 8186 7108 8188
rect 7164 8186 7188 8188
rect 7244 8186 7268 8188
rect 7324 8186 7330 8188
rect 7084 8134 7086 8186
rect 7266 8134 7268 8186
rect 7022 8132 7028 8134
rect 7084 8132 7108 8134
rect 7164 8132 7188 8134
rect 7244 8132 7268 8134
rect 7324 8132 7330 8134
rect 7022 8123 7330 8132
rect 9230 8188 9538 8197
rect 9230 8186 9236 8188
rect 9292 8186 9316 8188
rect 9372 8186 9396 8188
rect 9452 8186 9476 8188
rect 9532 8186 9538 8188
rect 9292 8134 9294 8186
rect 9474 8134 9476 8186
rect 9230 8132 9236 8134
rect 9292 8132 9316 8134
rect 9372 8132 9396 8134
rect 9452 8132 9476 8134
rect 9532 8132 9538 8134
rect 9230 8123 9538 8132
rect 1502 7644 1810 7653
rect 1502 7642 1508 7644
rect 1564 7642 1588 7644
rect 1644 7642 1668 7644
rect 1724 7642 1748 7644
rect 1804 7642 1810 7644
rect 1564 7590 1566 7642
rect 1746 7590 1748 7642
rect 1502 7588 1508 7590
rect 1564 7588 1588 7590
rect 1644 7588 1668 7590
rect 1724 7588 1748 7590
rect 1804 7588 1810 7590
rect 1502 7579 1810 7588
rect 3710 7644 4018 7653
rect 3710 7642 3716 7644
rect 3772 7642 3796 7644
rect 3852 7642 3876 7644
rect 3932 7642 3956 7644
rect 4012 7642 4018 7644
rect 3772 7590 3774 7642
rect 3954 7590 3956 7642
rect 3710 7588 3716 7590
rect 3772 7588 3796 7590
rect 3852 7588 3876 7590
rect 3932 7588 3956 7590
rect 4012 7588 4018 7590
rect 3710 7579 4018 7588
rect 5918 7644 6226 7653
rect 5918 7642 5924 7644
rect 5980 7642 6004 7644
rect 6060 7642 6084 7644
rect 6140 7642 6164 7644
rect 6220 7642 6226 7644
rect 5980 7590 5982 7642
rect 6162 7590 6164 7642
rect 5918 7588 5924 7590
rect 5980 7588 6004 7590
rect 6060 7588 6084 7590
rect 6140 7588 6164 7590
rect 6220 7588 6226 7590
rect 5918 7579 6226 7588
rect 8126 7644 8434 7653
rect 8126 7642 8132 7644
rect 8188 7642 8212 7644
rect 8268 7642 8292 7644
rect 8348 7642 8372 7644
rect 8428 7642 8434 7644
rect 8188 7590 8190 7642
rect 8370 7590 8372 7642
rect 8126 7588 8132 7590
rect 8188 7588 8212 7590
rect 8268 7588 8292 7590
rect 8348 7588 8372 7590
rect 8428 7588 8434 7590
rect 8126 7579 8434 7588
rect 2606 7100 2914 7109
rect 2606 7098 2612 7100
rect 2668 7098 2692 7100
rect 2748 7098 2772 7100
rect 2828 7098 2852 7100
rect 2908 7098 2914 7100
rect 2668 7046 2670 7098
rect 2850 7046 2852 7098
rect 2606 7044 2612 7046
rect 2668 7044 2692 7046
rect 2748 7044 2772 7046
rect 2828 7044 2852 7046
rect 2908 7044 2914 7046
rect 2606 7035 2914 7044
rect 4814 7100 5122 7109
rect 4814 7098 4820 7100
rect 4876 7098 4900 7100
rect 4956 7098 4980 7100
rect 5036 7098 5060 7100
rect 5116 7098 5122 7100
rect 4876 7046 4878 7098
rect 5058 7046 5060 7098
rect 4814 7044 4820 7046
rect 4876 7044 4900 7046
rect 4956 7044 4980 7046
rect 5036 7044 5060 7046
rect 5116 7044 5122 7046
rect 4814 7035 5122 7044
rect 7022 7100 7330 7109
rect 7022 7098 7028 7100
rect 7084 7098 7108 7100
rect 7164 7098 7188 7100
rect 7244 7098 7268 7100
rect 7324 7098 7330 7100
rect 7084 7046 7086 7098
rect 7266 7046 7268 7098
rect 7022 7044 7028 7046
rect 7084 7044 7108 7046
rect 7164 7044 7188 7046
rect 7244 7044 7268 7046
rect 7324 7044 7330 7046
rect 7022 7035 7330 7044
rect 9230 7100 9538 7109
rect 9230 7098 9236 7100
rect 9292 7098 9316 7100
rect 9372 7098 9396 7100
rect 9452 7098 9476 7100
rect 9532 7098 9538 7100
rect 9292 7046 9294 7098
rect 9474 7046 9476 7098
rect 9230 7044 9236 7046
rect 9292 7044 9316 7046
rect 9372 7044 9396 7046
rect 9452 7044 9476 7046
rect 9532 7044 9538 7046
rect 9230 7035 9538 7044
rect 1502 6556 1810 6565
rect 1502 6554 1508 6556
rect 1564 6554 1588 6556
rect 1644 6554 1668 6556
rect 1724 6554 1748 6556
rect 1804 6554 1810 6556
rect 1564 6502 1566 6554
rect 1746 6502 1748 6554
rect 1502 6500 1508 6502
rect 1564 6500 1588 6502
rect 1644 6500 1668 6502
rect 1724 6500 1748 6502
rect 1804 6500 1810 6502
rect 1502 6491 1810 6500
rect 3710 6556 4018 6565
rect 3710 6554 3716 6556
rect 3772 6554 3796 6556
rect 3852 6554 3876 6556
rect 3932 6554 3956 6556
rect 4012 6554 4018 6556
rect 3772 6502 3774 6554
rect 3954 6502 3956 6554
rect 3710 6500 3716 6502
rect 3772 6500 3796 6502
rect 3852 6500 3876 6502
rect 3932 6500 3956 6502
rect 4012 6500 4018 6502
rect 3710 6491 4018 6500
rect 5918 6556 6226 6565
rect 5918 6554 5924 6556
rect 5980 6554 6004 6556
rect 6060 6554 6084 6556
rect 6140 6554 6164 6556
rect 6220 6554 6226 6556
rect 5980 6502 5982 6554
rect 6162 6502 6164 6554
rect 5918 6500 5924 6502
rect 5980 6500 6004 6502
rect 6060 6500 6084 6502
rect 6140 6500 6164 6502
rect 6220 6500 6226 6502
rect 5918 6491 6226 6500
rect 8126 6556 8434 6565
rect 8126 6554 8132 6556
rect 8188 6554 8212 6556
rect 8268 6554 8292 6556
rect 8348 6554 8372 6556
rect 8428 6554 8434 6556
rect 8188 6502 8190 6554
rect 8370 6502 8372 6554
rect 8126 6500 8132 6502
rect 8188 6500 8212 6502
rect 8268 6500 8292 6502
rect 8348 6500 8372 6502
rect 8428 6500 8434 6502
rect 8126 6491 8434 6500
rect 2606 6012 2914 6021
rect 2606 6010 2612 6012
rect 2668 6010 2692 6012
rect 2748 6010 2772 6012
rect 2828 6010 2852 6012
rect 2908 6010 2914 6012
rect 2668 5958 2670 6010
rect 2850 5958 2852 6010
rect 2606 5956 2612 5958
rect 2668 5956 2692 5958
rect 2748 5956 2772 5958
rect 2828 5956 2852 5958
rect 2908 5956 2914 5958
rect 2606 5947 2914 5956
rect 4814 6012 5122 6021
rect 4814 6010 4820 6012
rect 4876 6010 4900 6012
rect 4956 6010 4980 6012
rect 5036 6010 5060 6012
rect 5116 6010 5122 6012
rect 4876 5958 4878 6010
rect 5058 5958 5060 6010
rect 4814 5956 4820 5958
rect 4876 5956 4900 5958
rect 4956 5956 4980 5958
rect 5036 5956 5060 5958
rect 5116 5956 5122 5958
rect 4814 5947 5122 5956
rect 7022 6012 7330 6021
rect 7022 6010 7028 6012
rect 7084 6010 7108 6012
rect 7164 6010 7188 6012
rect 7244 6010 7268 6012
rect 7324 6010 7330 6012
rect 7084 5958 7086 6010
rect 7266 5958 7268 6010
rect 7022 5956 7028 5958
rect 7084 5956 7108 5958
rect 7164 5956 7188 5958
rect 7244 5956 7268 5958
rect 7324 5956 7330 5958
rect 7022 5947 7330 5956
rect 9230 6012 9538 6021
rect 9230 6010 9236 6012
rect 9292 6010 9316 6012
rect 9372 6010 9396 6012
rect 9452 6010 9476 6012
rect 9532 6010 9538 6012
rect 9292 5958 9294 6010
rect 9474 5958 9476 6010
rect 9230 5956 9236 5958
rect 9292 5956 9316 5958
rect 9372 5956 9396 5958
rect 9452 5956 9476 5958
rect 9532 5956 9538 5958
rect 9230 5947 9538 5956
rect 1502 5468 1810 5477
rect 1502 5466 1508 5468
rect 1564 5466 1588 5468
rect 1644 5466 1668 5468
rect 1724 5466 1748 5468
rect 1804 5466 1810 5468
rect 1564 5414 1566 5466
rect 1746 5414 1748 5466
rect 1502 5412 1508 5414
rect 1564 5412 1588 5414
rect 1644 5412 1668 5414
rect 1724 5412 1748 5414
rect 1804 5412 1810 5414
rect 1502 5403 1810 5412
rect 3710 5468 4018 5477
rect 3710 5466 3716 5468
rect 3772 5466 3796 5468
rect 3852 5466 3876 5468
rect 3932 5466 3956 5468
rect 4012 5466 4018 5468
rect 3772 5414 3774 5466
rect 3954 5414 3956 5466
rect 3710 5412 3716 5414
rect 3772 5412 3796 5414
rect 3852 5412 3876 5414
rect 3932 5412 3956 5414
rect 4012 5412 4018 5414
rect 3710 5403 4018 5412
rect 5918 5468 6226 5477
rect 5918 5466 5924 5468
rect 5980 5466 6004 5468
rect 6060 5466 6084 5468
rect 6140 5466 6164 5468
rect 6220 5466 6226 5468
rect 5980 5414 5982 5466
rect 6162 5414 6164 5466
rect 5918 5412 5924 5414
rect 5980 5412 6004 5414
rect 6060 5412 6084 5414
rect 6140 5412 6164 5414
rect 6220 5412 6226 5414
rect 5918 5403 6226 5412
rect 8126 5468 8434 5477
rect 8126 5466 8132 5468
rect 8188 5466 8212 5468
rect 8268 5466 8292 5468
rect 8348 5466 8372 5468
rect 8428 5466 8434 5468
rect 8188 5414 8190 5466
rect 8370 5414 8372 5466
rect 8126 5412 8132 5414
rect 8188 5412 8212 5414
rect 8268 5412 8292 5414
rect 8348 5412 8372 5414
rect 8428 5412 8434 5414
rect 8126 5403 8434 5412
rect 2606 4924 2914 4933
rect 2606 4922 2612 4924
rect 2668 4922 2692 4924
rect 2748 4922 2772 4924
rect 2828 4922 2852 4924
rect 2908 4922 2914 4924
rect 2668 4870 2670 4922
rect 2850 4870 2852 4922
rect 2606 4868 2612 4870
rect 2668 4868 2692 4870
rect 2748 4868 2772 4870
rect 2828 4868 2852 4870
rect 2908 4868 2914 4870
rect 2606 4859 2914 4868
rect 4814 4924 5122 4933
rect 4814 4922 4820 4924
rect 4876 4922 4900 4924
rect 4956 4922 4980 4924
rect 5036 4922 5060 4924
rect 5116 4922 5122 4924
rect 4876 4870 4878 4922
rect 5058 4870 5060 4922
rect 4814 4868 4820 4870
rect 4876 4868 4900 4870
rect 4956 4868 4980 4870
rect 5036 4868 5060 4870
rect 5116 4868 5122 4870
rect 4814 4859 5122 4868
rect 7022 4924 7330 4933
rect 7022 4922 7028 4924
rect 7084 4922 7108 4924
rect 7164 4922 7188 4924
rect 7244 4922 7268 4924
rect 7324 4922 7330 4924
rect 7084 4870 7086 4922
rect 7266 4870 7268 4922
rect 7022 4868 7028 4870
rect 7084 4868 7108 4870
rect 7164 4868 7188 4870
rect 7244 4868 7268 4870
rect 7324 4868 7330 4870
rect 7022 4859 7330 4868
rect 9230 4924 9538 4933
rect 9230 4922 9236 4924
rect 9292 4922 9316 4924
rect 9372 4922 9396 4924
rect 9452 4922 9476 4924
rect 9532 4922 9538 4924
rect 9292 4870 9294 4922
rect 9474 4870 9476 4922
rect 9230 4868 9236 4870
rect 9292 4868 9316 4870
rect 9372 4868 9396 4870
rect 9452 4868 9476 4870
rect 9532 4868 9538 4870
rect 9230 4859 9538 4868
rect 1502 4380 1810 4389
rect 1502 4378 1508 4380
rect 1564 4378 1588 4380
rect 1644 4378 1668 4380
rect 1724 4378 1748 4380
rect 1804 4378 1810 4380
rect 1564 4326 1566 4378
rect 1746 4326 1748 4378
rect 1502 4324 1508 4326
rect 1564 4324 1588 4326
rect 1644 4324 1668 4326
rect 1724 4324 1748 4326
rect 1804 4324 1810 4326
rect 1502 4315 1810 4324
rect 3710 4380 4018 4389
rect 3710 4378 3716 4380
rect 3772 4378 3796 4380
rect 3852 4378 3876 4380
rect 3932 4378 3956 4380
rect 4012 4378 4018 4380
rect 3772 4326 3774 4378
rect 3954 4326 3956 4378
rect 3710 4324 3716 4326
rect 3772 4324 3796 4326
rect 3852 4324 3876 4326
rect 3932 4324 3956 4326
rect 4012 4324 4018 4326
rect 3710 4315 4018 4324
rect 5918 4380 6226 4389
rect 5918 4378 5924 4380
rect 5980 4378 6004 4380
rect 6060 4378 6084 4380
rect 6140 4378 6164 4380
rect 6220 4378 6226 4380
rect 5980 4326 5982 4378
rect 6162 4326 6164 4378
rect 5918 4324 5924 4326
rect 5980 4324 6004 4326
rect 6060 4324 6084 4326
rect 6140 4324 6164 4326
rect 6220 4324 6226 4326
rect 5918 4315 6226 4324
rect 8126 4380 8434 4389
rect 8126 4378 8132 4380
rect 8188 4378 8212 4380
rect 8268 4378 8292 4380
rect 8348 4378 8372 4380
rect 8428 4378 8434 4380
rect 8188 4326 8190 4378
rect 8370 4326 8372 4378
rect 8126 4324 8132 4326
rect 8188 4324 8212 4326
rect 8268 4324 8292 4326
rect 8348 4324 8372 4326
rect 8428 4324 8434 4326
rect 8126 4315 8434 4324
rect 2606 3836 2914 3845
rect 2606 3834 2612 3836
rect 2668 3834 2692 3836
rect 2748 3834 2772 3836
rect 2828 3834 2852 3836
rect 2908 3834 2914 3836
rect 2668 3782 2670 3834
rect 2850 3782 2852 3834
rect 2606 3780 2612 3782
rect 2668 3780 2692 3782
rect 2748 3780 2772 3782
rect 2828 3780 2852 3782
rect 2908 3780 2914 3782
rect 2606 3771 2914 3780
rect 4814 3836 5122 3845
rect 4814 3834 4820 3836
rect 4876 3834 4900 3836
rect 4956 3834 4980 3836
rect 5036 3834 5060 3836
rect 5116 3834 5122 3836
rect 4876 3782 4878 3834
rect 5058 3782 5060 3834
rect 4814 3780 4820 3782
rect 4876 3780 4900 3782
rect 4956 3780 4980 3782
rect 5036 3780 5060 3782
rect 5116 3780 5122 3782
rect 4814 3771 5122 3780
rect 7022 3836 7330 3845
rect 7022 3834 7028 3836
rect 7084 3834 7108 3836
rect 7164 3834 7188 3836
rect 7244 3834 7268 3836
rect 7324 3834 7330 3836
rect 7084 3782 7086 3834
rect 7266 3782 7268 3834
rect 7022 3780 7028 3782
rect 7084 3780 7108 3782
rect 7164 3780 7188 3782
rect 7244 3780 7268 3782
rect 7324 3780 7330 3782
rect 7022 3771 7330 3780
rect 9230 3836 9538 3845
rect 9230 3834 9236 3836
rect 9292 3834 9316 3836
rect 9372 3834 9396 3836
rect 9452 3834 9476 3836
rect 9532 3834 9538 3836
rect 9292 3782 9294 3834
rect 9474 3782 9476 3834
rect 9230 3780 9236 3782
rect 9292 3780 9316 3782
rect 9372 3780 9396 3782
rect 9452 3780 9476 3782
rect 9532 3780 9538 3782
rect 9230 3771 9538 3780
rect 1502 3292 1810 3301
rect 1502 3290 1508 3292
rect 1564 3290 1588 3292
rect 1644 3290 1668 3292
rect 1724 3290 1748 3292
rect 1804 3290 1810 3292
rect 1564 3238 1566 3290
rect 1746 3238 1748 3290
rect 1502 3236 1508 3238
rect 1564 3236 1588 3238
rect 1644 3236 1668 3238
rect 1724 3236 1748 3238
rect 1804 3236 1810 3238
rect 1502 3227 1810 3236
rect 3710 3292 4018 3301
rect 3710 3290 3716 3292
rect 3772 3290 3796 3292
rect 3852 3290 3876 3292
rect 3932 3290 3956 3292
rect 4012 3290 4018 3292
rect 3772 3238 3774 3290
rect 3954 3238 3956 3290
rect 3710 3236 3716 3238
rect 3772 3236 3796 3238
rect 3852 3236 3876 3238
rect 3932 3236 3956 3238
rect 4012 3236 4018 3238
rect 3710 3227 4018 3236
rect 5918 3292 6226 3301
rect 5918 3290 5924 3292
rect 5980 3290 6004 3292
rect 6060 3290 6084 3292
rect 6140 3290 6164 3292
rect 6220 3290 6226 3292
rect 5980 3238 5982 3290
rect 6162 3238 6164 3290
rect 5918 3236 5924 3238
rect 5980 3236 6004 3238
rect 6060 3236 6084 3238
rect 6140 3236 6164 3238
rect 6220 3236 6226 3238
rect 5918 3227 6226 3236
rect 8126 3292 8434 3301
rect 8126 3290 8132 3292
rect 8188 3290 8212 3292
rect 8268 3290 8292 3292
rect 8348 3290 8372 3292
rect 8428 3290 8434 3292
rect 8188 3238 8190 3290
rect 8370 3238 8372 3290
rect 8126 3236 8132 3238
rect 8188 3236 8212 3238
rect 8268 3236 8292 3238
rect 8348 3236 8372 3238
rect 8428 3236 8434 3238
rect 8126 3227 8434 3236
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 2606 2748 2914 2757
rect 2606 2746 2612 2748
rect 2668 2746 2692 2748
rect 2748 2746 2772 2748
rect 2828 2746 2852 2748
rect 2908 2746 2914 2748
rect 2668 2694 2670 2746
rect 2850 2694 2852 2746
rect 2606 2692 2612 2694
rect 2668 2692 2692 2694
rect 2748 2692 2772 2694
rect 2828 2692 2852 2694
rect 2908 2692 2914 2694
rect 2606 2683 2914 2692
rect 4172 2650 4200 2926
rect 4814 2748 5122 2757
rect 4814 2746 4820 2748
rect 4876 2746 4900 2748
rect 4956 2746 4980 2748
rect 5036 2746 5060 2748
rect 5116 2746 5122 2748
rect 4876 2694 4878 2746
rect 5058 2694 5060 2746
rect 4814 2692 4820 2694
rect 4876 2692 4900 2694
rect 4956 2692 4980 2694
rect 5036 2692 5060 2694
rect 5116 2692 5122 2694
rect 4814 2683 5122 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 1502 2204 1810 2213
rect 1502 2202 1508 2204
rect 1564 2202 1588 2204
rect 1644 2202 1668 2204
rect 1724 2202 1748 2204
rect 1804 2202 1810 2204
rect 1564 2150 1566 2202
rect 1746 2150 1748 2202
rect 1502 2148 1508 2150
rect 1564 2148 1588 2150
rect 1644 2148 1668 2150
rect 1724 2148 1748 2150
rect 1804 2148 1810 2150
rect 1502 2139 1810 2148
rect 3710 2204 4018 2213
rect 3710 2202 3716 2204
rect 3772 2202 3796 2204
rect 3852 2202 3876 2204
rect 3932 2202 3956 2204
rect 4012 2202 4018 2204
rect 3772 2150 3774 2202
rect 3954 2150 3956 2202
rect 3710 2148 3716 2150
rect 3772 2148 3796 2150
rect 3852 2148 3876 2150
rect 3932 2148 3956 2150
rect 4012 2148 4018 2150
rect 3710 2139 4018 2148
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 2516 1562 2544 1838
rect 3424 1828 3476 1834
rect 3424 1770 3476 1776
rect 3056 1760 3108 1766
rect 3056 1702 3108 1708
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 2606 1660 2914 1669
rect 2606 1658 2612 1660
rect 2668 1658 2692 1660
rect 2748 1658 2772 1660
rect 2828 1658 2852 1660
rect 2908 1658 2914 1660
rect 2668 1606 2670 1658
rect 2850 1606 2852 1658
rect 2606 1604 2612 1606
rect 2668 1604 2692 1606
rect 2748 1604 2772 1606
rect 2828 1604 2852 1606
rect 2908 1604 2914 1606
rect 2606 1595 2914 1604
rect 2504 1556 2556 1562
rect 2504 1498 2556 1504
rect 3068 1426 3096 1702
rect 3252 1494 3280 1702
rect 3240 1488 3292 1494
rect 3240 1430 3292 1436
rect 2320 1420 2372 1426
rect 2320 1362 2372 1368
rect 3056 1420 3108 1426
rect 3056 1362 3108 1368
rect 1308 1352 1360 1358
rect 1308 1294 1360 1300
rect 1320 678 1348 1294
rect 1502 1116 1810 1125
rect 1502 1114 1508 1116
rect 1564 1114 1588 1116
rect 1644 1114 1668 1116
rect 1724 1114 1748 1116
rect 1804 1114 1810 1116
rect 1564 1062 1566 1114
rect 1746 1062 1748 1114
rect 1502 1060 1508 1062
rect 1564 1060 1588 1062
rect 1644 1060 1668 1062
rect 1724 1060 1748 1062
rect 1804 1060 1810 1062
rect 1502 1051 1810 1060
rect 2332 1018 2360 1362
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 2320 1012 2372 1018
rect 2320 954 2372 960
rect 2516 814 2544 1158
rect 3436 1018 3464 1770
rect 3804 1222 3832 1838
rect 4172 1426 4200 2586
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4252 2032 4304 2038
rect 4252 1974 4304 1980
rect 4160 1420 4212 1426
rect 4160 1362 4212 1368
rect 3792 1216 3844 1222
rect 3792 1158 3844 1164
rect 3710 1116 4018 1125
rect 3710 1114 3716 1116
rect 3772 1114 3796 1116
rect 3852 1114 3876 1116
rect 3932 1114 3956 1116
rect 4012 1114 4018 1116
rect 3772 1062 3774 1114
rect 3954 1062 3956 1114
rect 3710 1060 3716 1062
rect 3772 1060 3796 1062
rect 3852 1060 3876 1062
rect 3932 1060 3956 1062
rect 4012 1060 4018 1062
rect 3710 1051 4018 1060
rect 3424 1012 3476 1018
rect 3424 954 3476 960
rect 4172 882 4200 1362
rect 4160 876 4212 882
rect 4160 818 4212 824
rect 4264 814 4292 1974
rect 4448 1766 4476 2450
rect 4712 1896 4764 1902
rect 4712 1838 4764 1844
rect 4436 1760 4488 1766
rect 4436 1702 4488 1708
rect 4724 1562 4752 1838
rect 4814 1660 5122 1669
rect 4814 1658 4820 1660
rect 4876 1658 4900 1660
rect 4956 1658 4980 1660
rect 5036 1658 5060 1660
rect 5116 1658 5122 1660
rect 4876 1606 4878 1658
rect 5058 1606 5060 1658
rect 4814 1604 4820 1606
rect 4876 1604 4900 1606
rect 4956 1604 4980 1606
rect 5036 1604 5060 1606
rect 5116 1604 5122 1606
rect 4814 1595 5122 1604
rect 4712 1556 4764 1562
rect 4712 1498 4764 1504
rect 4896 1352 4948 1358
rect 4896 1294 4948 1300
rect 4436 1216 4488 1222
rect 4436 1158 4488 1164
rect 2504 808 2556 814
rect 2504 750 2556 756
rect 4252 808 4304 814
rect 4252 750 4304 756
rect 848 672 900 678
rect 848 614 900 620
rect 1308 672 1360 678
rect 1308 614 1360 620
rect 860 400 888 614
rect 2516 400 2544 750
rect 4448 678 4476 1158
rect 4908 678 4936 1294
rect 5184 1018 5212 2926
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5368 1222 5396 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 5356 1216 5408 1222
rect 5356 1158 5408 1164
rect 5460 1018 5488 2314
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5172 1012 5224 1018
rect 5172 954 5224 960
rect 5448 1012 5500 1018
rect 5448 954 5500 960
rect 5552 814 5580 2246
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5644 950 5672 1362
rect 5828 1358 5856 2790
rect 7022 2748 7330 2757
rect 7022 2746 7028 2748
rect 7084 2746 7108 2748
rect 7164 2746 7188 2748
rect 7244 2746 7268 2748
rect 7324 2746 7330 2748
rect 7084 2694 7086 2746
rect 7266 2694 7268 2746
rect 7022 2692 7028 2694
rect 7084 2692 7108 2694
rect 7164 2692 7188 2694
rect 7244 2692 7268 2694
rect 7324 2692 7330 2694
rect 7022 2683 7330 2692
rect 9230 2748 9538 2757
rect 9230 2746 9236 2748
rect 9292 2746 9316 2748
rect 9372 2746 9396 2748
rect 9452 2746 9476 2748
rect 9532 2746 9538 2748
rect 9292 2694 9294 2746
rect 9474 2694 9476 2746
rect 9230 2692 9236 2694
rect 9292 2692 9316 2694
rect 9372 2692 9396 2694
rect 9452 2692 9476 2694
rect 9532 2692 9538 2694
rect 9230 2683 9538 2692
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 5918 2204 6226 2213
rect 5918 2202 5924 2204
rect 5980 2202 6004 2204
rect 6060 2202 6084 2204
rect 6140 2202 6164 2204
rect 6220 2202 6226 2204
rect 5980 2150 5982 2202
rect 6162 2150 6164 2202
rect 5918 2148 5924 2150
rect 5980 2148 6004 2150
rect 6060 2148 6084 2150
rect 6140 2148 6164 2150
rect 6220 2148 6226 2150
rect 5918 2139 6226 2148
rect 6276 1556 6328 1562
rect 6276 1498 6328 1504
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 5632 944 5684 950
rect 5632 886 5684 892
rect 5540 808 5592 814
rect 5540 750 5592 756
rect 2964 672 3016 678
rect 2964 614 3016 620
rect 4436 672 4488 678
rect 4436 614 4488 620
rect 4528 672 4580 678
rect 4528 614 4580 620
rect 4896 672 4948 678
rect 4896 614 4948 620
rect 2606 572 2914 581
rect 2606 570 2612 572
rect 2668 570 2692 572
rect 2748 570 2772 572
rect 2828 570 2852 572
rect 2908 570 2914 572
rect 2668 518 2670 570
rect 2850 518 2852 570
rect 2606 516 2612 518
rect 2668 516 2692 518
rect 2748 516 2772 518
rect 2828 516 2852 518
rect 2908 516 2914 518
rect 2606 507 2914 516
rect 2976 474 3004 614
rect 2964 468 3016 474
rect 2964 410 3016 416
rect 4172 462 4292 490
rect 4172 400 4200 462
rect 846 0 902 400
rect 2502 0 2558 400
rect 4158 0 4214 400
rect 4264 354 4292 462
rect 4540 354 4568 614
rect 4814 572 5122 581
rect 4814 570 4820 572
rect 4876 570 4900 572
rect 4956 570 4980 572
rect 5036 570 5060 572
rect 5116 570 5122 572
rect 4876 518 4878 570
rect 5058 518 5060 570
rect 4814 516 4820 518
rect 4876 516 4900 518
rect 4956 516 4980 518
rect 5036 516 5060 518
rect 5116 516 5122 518
rect 4814 507 5122 516
rect 5736 474 5764 1294
rect 5828 882 5856 1294
rect 5918 1116 6226 1125
rect 5918 1114 5924 1116
rect 5980 1114 6004 1116
rect 6060 1114 6084 1116
rect 6140 1114 6164 1116
rect 6220 1114 6226 1116
rect 5980 1062 5982 1114
rect 6162 1062 6164 1114
rect 5918 1060 5924 1062
rect 5980 1060 6004 1062
rect 6060 1060 6084 1062
rect 6140 1060 6164 1062
rect 6220 1060 6226 1062
rect 5918 1051 6226 1060
rect 5816 876 5868 882
rect 5816 818 5868 824
rect 5724 468 5776 474
rect 5724 410 5776 416
rect 5828 400 5856 818
rect 6288 746 6316 1498
rect 6380 1426 6408 2246
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 6460 1760 6512 1766
rect 6460 1702 6512 1708
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 6380 814 6408 1362
rect 6472 814 6500 1702
rect 6748 1426 6776 1838
rect 7472 1828 7524 1834
rect 7472 1770 7524 1776
rect 7380 1760 7432 1766
rect 7380 1702 7432 1708
rect 7022 1660 7330 1669
rect 7022 1658 7028 1660
rect 7084 1658 7108 1660
rect 7164 1658 7188 1660
rect 7244 1658 7268 1660
rect 7324 1658 7330 1660
rect 7084 1606 7086 1658
rect 7266 1606 7268 1658
rect 7022 1604 7028 1606
rect 7084 1604 7108 1606
rect 7164 1604 7188 1606
rect 7244 1604 7268 1606
rect 7324 1604 7330 1606
rect 7022 1595 7330 1604
rect 7392 1494 7420 1702
rect 7380 1488 7432 1494
rect 7380 1430 7432 1436
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 6748 950 6776 1362
rect 6736 944 6788 950
rect 6736 886 6788 892
rect 6368 808 6420 814
rect 6368 750 6420 756
rect 6460 808 6512 814
rect 6460 750 6512 756
rect 6276 740 6328 746
rect 6276 682 6328 688
rect 7022 572 7330 581
rect 7022 570 7028 572
rect 7084 570 7108 572
rect 7164 570 7188 572
rect 7244 570 7268 572
rect 7324 570 7330 572
rect 7084 518 7086 570
rect 7266 518 7268 570
rect 7022 516 7028 518
rect 7084 516 7108 518
rect 7164 516 7188 518
rect 7244 516 7268 518
rect 7324 516 7330 518
rect 7022 507 7330 516
rect 7484 400 7512 1770
rect 7944 1562 7972 2382
rect 8126 2204 8434 2213
rect 8126 2202 8132 2204
rect 8188 2202 8212 2204
rect 8268 2202 8292 2204
rect 8348 2202 8372 2204
rect 8428 2202 8434 2204
rect 8188 2150 8190 2202
rect 8370 2150 8372 2202
rect 8126 2148 8132 2150
rect 8188 2148 8212 2150
rect 8268 2148 8292 2150
rect 8348 2148 8372 2150
rect 8428 2148 8434 2150
rect 8126 2139 8434 2148
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 7944 1018 7972 1498
rect 8588 1358 8616 2382
rect 8944 1896 8996 1902
rect 8944 1838 8996 1844
rect 8852 1420 8904 1426
rect 8852 1362 8904 1368
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 8126 1116 8434 1125
rect 8126 1114 8132 1116
rect 8188 1114 8212 1116
rect 8268 1114 8292 1116
rect 8348 1114 8372 1116
rect 8428 1114 8434 1116
rect 8188 1062 8190 1114
rect 8370 1062 8372 1114
rect 8126 1060 8132 1062
rect 8188 1060 8212 1062
rect 8268 1060 8292 1062
rect 8348 1060 8372 1062
rect 8428 1060 8434 1062
rect 8126 1051 8434 1060
rect 8864 1018 8892 1362
rect 8956 1222 8984 1838
rect 9230 1660 9538 1669
rect 9230 1658 9236 1660
rect 9292 1658 9316 1660
rect 9372 1658 9396 1660
rect 9452 1658 9476 1660
rect 9532 1658 9538 1660
rect 9292 1606 9294 1658
rect 9474 1606 9476 1658
rect 9230 1604 9236 1606
rect 9292 1604 9316 1606
rect 9372 1604 9396 1606
rect 9452 1604 9476 1606
rect 9532 1604 9538 1606
rect 9230 1595 9538 1604
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 7932 1012 7984 1018
rect 7932 954 7984 960
rect 8852 1012 8904 1018
rect 8852 954 8904 960
rect 9128 808 9180 814
rect 9128 750 9180 756
rect 9140 400 9168 750
rect 9230 572 9538 581
rect 9230 570 9236 572
rect 9292 570 9316 572
rect 9372 570 9396 572
rect 9452 570 9476 572
rect 9532 570 9538 572
rect 9292 518 9294 570
rect 9474 518 9476 570
rect 9230 516 9236 518
rect 9292 516 9316 518
rect 9372 516 9396 518
rect 9452 516 9476 518
rect 9532 516 9538 518
rect 9230 507 9538 516
rect 4264 326 4568 354
rect 5814 0 5870 400
rect 7470 0 7526 400
rect 9126 0 9182 400
<< via2 >>
rect 2612 9274 2668 9276
rect 2692 9274 2748 9276
rect 2772 9274 2828 9276
rect 2852 9274 2908 9276
rect 2612 9222 2658 9274
rect 2658 9222 2668 9274
rect 2692 9222 2722 9274
rect 2722 9222 2734 9274
rect 2734 9222 2748 9274
rect 2772 9222 2786 9274
rect 2786 9222 2798 9274
rect 2798 9222 2828 9274
rect 2852 9222 2862 9274
rect 2862 9222 2908 9274
rect 2612 9220 2668 9222
rect 2692 9220 2748 9222
rect 2772 9220 2828 9222
rect 2852 9220 2908 9222
rect 4820 9274 4876 9276
rect 4900 9274 4956 9276
rect 4980 9274 5036 9276
rect 5060 9274 5116 9276
rect 4820 9222 4866 9274
rect 4866 9222 4876 9274
rect 4900 9222 4930 9274
rect 4930 9222 4942 9274
rect 4942 9222 4956 9274
rect 4980 9222 4994 9274
rect 4994 9222 5006 9274
rect 5006 9222 5036 9274
rect 5060 9222 5070 9274
rect 5070 9222 5116 9274
rect 4820 9220 4876 9222
rect 4900 9220 4956 9222
rect 4980 9220 5036 9222
rect 5060 9220 5116 9222
rect 7028 9274 7084 9276
rect 7108 9274 7164 9276
rect 7188 9274 7244 9276
rect 7268 9274 7324 9276
rect 7028 9222 7074 9274
rect 7074 9222 7084 9274
rect 7108 9222 7138 9274
rect 7138 9222 7150 9274
rect 7150 9222 7164 9274
rect 7188 9222 7202 9274
rect 7202 9222 7214 9274
rect 7214 9222 7244 9274
rect 7268 9222 7278 9274
rect 7278 9222 7324 9274
rect 7028 9220 7084 9222
rect 7108 9220 7164 9222
rect 7188 9220 7244 9222
rect 7268 9220 7324 9222
rect 9236 9274 9292 9276
rect 9316 9274 9372 9276
rect 9396 9274 9452 9276
rect 9476 9274 9532 9276
rect 9236 9222 9282 9274
rect 9282 9222 9292 9274
rect 9316 9222 9346 9274
rect 9346 9222 9358 9274
rect 9358 9222 9372 9274
rect 9396 9222 9410 9274
rect 9410 9222 9422 9274
rect 9422 9222 9452 9274
rect 9476 9222 9486 9274
rect 9486 9222 9532 9274
rect 9236 9220 9292 9222
rect 9316 9220 9372 9222
rect 9396 9220 9452 9222
rect 9476 9220 9532 9222
rect 1508 8730 1564 8732
rect 1588 8730 1644 8732
rect 1668 8730 1724 8732
rect 1748 8730 1804 8732
rect 1508 8678 1554 8730
rect 1554 8678 1564 8730
rect 1588 8678 1618 8730
rect 1618 8678 1630 8730
rect 1630 8678 1644 8730
rect 1668 8678 1682 8730
rect 1682 8678 1694 8730
rect 1694 8678 1724 8730
rect 1748 8678 1758 8730
rect 1758 8678 1804 8730
rect 1508 8676 1564 8678
rect 1588 8676 1644 8678
rect 1668 8676 1724 8678
rect 1748 8676 1804 8678
rect 3716 8730 3772 8732
rect 3796 8730 3852 8732
rect 3876 8730 3932 8732
rect 3956 8730 4012 8732
rect 3716 8678 3762 8730
rect 3762 8678 3772 8730
rect 3796 8678 3826 8730
rect 3826 8678 3838 8730
rect 3838 8678 3852 8730
rect 3876 8678 3890 8730
rect 3890 8678 3902 8730
rect 3902 8678 3932 8730
rect 3956 8678 3966 8730
rect 3966 8678 4012 8730
rect 3716 8676 3772 8678
rect 3796 8676 3852 8678
rect 3876 8676 3932 8678
rect 3956 8676 4012 8678
rect 5924 8730 5980 8732
rect 6004 8730 6060 8732
rect 6084 8730 6140 8732
rect 6164 8730 6220 8732
rect 5924 8678 5970 8730
rect 5970 8678 5980 8730
rect 6004 8678 6034 8730
rect 6034 8678 6046 8730
rect 6046 8678 6060 8730
rect 6084 8678 6098 8730
rect 6098 8678 6110 8730
rect 6110 8678 6140 8730
rect 6164 8678 6174 8730
rect 6174 8678 6220 8730
rect 5924 8676 5980 8678
rect 6004 8676 6060 8678
rect 6084 8676 6140 8678
rect 6164 8676 6220 8678
rect 8132 8730 8188 8732
rect 8212 8730 8268 8732
rect 8292 8730 8348 8732
rect 8372 8730 8428 8732
rect 8132 8678 8178 8730
rect 8178 8678 8188 8730
rect 8212 8678 8242 8730
rect 8242 8678 8254 8730
rect 8254 8678 8268 8730
rect 8292 8678 8306 8730
rect 8306 8678 8318 8730
rect 8318 8678 8348 8730
rect 8372 8678 8382 8730
rect 8382 8678 8428 8730
rect 8132 8676 8188 8678
rect 8212 8676 8268 8678
rect 8292 8676 8348 8678
rect 8372 8676 8428 8678
rect 2612 8186 2668 8188
rect 2692 8186 2748 8188
rect 2772 8186 2828 8188
rect 2852 8186 2908 8188
rect 2612 8134 2658 8186
rect 2658 8134 2668 8186
rect 2692 8134 2722 8186
rect 2722 8134 2734 8186
rect 2734 8134 2748 8186
rect 2772 8134 2786 8186
rect 2786 8134 2798 8186
rect 2798 8134 2828 8186
rect 2852 8134 2862 8186
rect 2862 8134 2908 8186
rect 2612 8132 2668 8134
rect 2692 8132 2748 8134
rect 2772 8132 2828 8134
rect 2852 8132 2908 8134
rect 4820 8186 4876 8188
rect 4900 8186 4956 8188
rect 4980 8186 5036 8188
rect 5060 8186 5116 8188
rect 4820 8134 4866 8186
rect 4866 8134 4876 8186
rect 4900 8134 4930 8186
rect 4930 8134 4942 8186
rect 4942 8134 4956 8186
rect 4980 8134 4994 8186
rect 4994 8134 5006 8186
rect 5006 8134 5036 8186
rect 5060 8134 5070 8186
rect 5070 8134 5116 8186
rect 4820 8132 4876 8134
rect 4900 8132 4956 8134
rect 4980 8132 5036 8134
rect 5060 8132 5116 8134
rect 7028 8186 7084 8188
rect 7108 8186 7164 8188
rect 7188 8186 7244 8188
rect 7268 8186 7324 8188
rect 7028 8134 7074 8186
rect 7074 8134 7084 8186
rect 7108 8134 7138 8186
rect 7138 8134 7150 8186
rect 7150 8134 7164 8186
rect 7188 8134 7202 8186
rect 7202 8134 7214 8186
rect 7214 8134 7244 8186
rect 7268 8134 7278 8186
rect 7278 8134 7324 8186
rect 7028 8132 7084 8134
rect 7108 8132 7164 8134
rect 7188 8132 7244 8134
rect 7268 8132 7324 8134
rect 9236 8186 9292 8188
rect 9316 8186 9372 8188
rect 9396 8186 9452 8188
rect 9476 8186 9532 8188
rect 9236 8134 9282 8186
rect 9282 8134 9292 8186
rect 9316 8134 9346 8186
rect 9346 8134 9358 8186
rect 9358 8134 9372 8186
rect 9396 8134 9410 8186
rect 9410 8134 9422 8186
rect 9422 8134 9452 8186
rect 9476 8134 9486 8186
rect 9486 8134 9532 8186
rect 9236 8132 9292 8134
rect 9316 8132 9372 8134
rect 9396 8132 9452 8134
rect 9476 8132 9532 8134
rect 1508 7642 1564 7644
rect 1588 7642 1644 7644
rect 1668 7642 1724 7644
rect 1748 7642 1804 7644
rect 1508 7590 1554 7642
rect 1554 7590 1564 7642
rect 1588 7590 1618 7642
rect 1618 7590 1630 7642
rect 1630 7590 1644 7642
rect 1668 7590 1682 7642
rect 1682 7590 1694 7642
rect 1694 7590 1724 7642
rect 1748 7590 1758 7642
rect 1758 7590 1804 7642
rect 1508 7588 1564 7590
rect 1588 7588 1644 7590
rect 1668 7588 1724 7590
rect 1748 7588 1804 7590
rect 3716 7642 3772 7644
rect 3796 7642 3852 7644
rect 3876 7642 3932 7644
rect 3956 7642 4012 7644
rect 3716 7590 3762 7642
rect 3762 7590 3772 7642
rect 3796 7590 3826 7642
rect 3826 7590 3838 7642
rect 3838 7590 3852 7642
rect 3876 7590 3890 7642
rect 3890 7590 3902 7642
rect 3902 7590 3932 7642
rect 3956 7590 3966 7642
rect 3966 7590 4012 7642
rect 3716 7588 3772 7590
rect 3796 7588 3852 7590
rect 3876 7588 3932 7590
rect 3956 7588 4012 7590
rect 5924 7642 5980 7644
rect 6004 7642 6060 7644
rect 6084 7642 6140 7644
rect 6164 7642 6220 7644
rect 5924 7590 5970 7642
rect 5970 7590 5980 7642
rect 6004 7590 6034 7642
rect 6034 7590 6046 7642
rect 6046 7590 6060 7642
rect 6084 7590 6098 7642
rect 6098 7590 6110 7642
rect 6110 7590 6140 7642
rect 6164 7590 6174 7642
rect 6174 7590 6220 7642
rect 5924 7588 5980 7590
rect 6004 7588 6060 7590
rect 6084 7588 6140 7590
rect 6164 7588 6220 7590
rect 8132 7642 8188 7644
rect 8212 7642 8268 7644
rect 8292 7642 8348 7644
rect 8372 7642 8428 7644
rect 8132 7590 8178 7642
rect 8178 7590 8188 7642
rect 8212 7590 8242 7642
rect 8242 7590 8254 7642
rect 8254 7590 8268 7642
rect 8292 7590 8306 7642
rect 8306 7590 8318 7642
rect 8318 7590 8348 7642
rect 8372 7590 8382 7642
rect 8382 7590 8428 7642
rect 8132 7588 8188 7590
rect 8212 7588 8268 7590
rect 8292 7588 8348 7590
rect 8372 7588 8428 7590
rect 2612 7098 2668 7100
rect 2692 7098 2748 7100
rect 2772 7098 2828 7100
rect 2852 7098 2908 7100
rect 2612 7046 2658 7098
rect 2658 7046 2668 7098
rect 2692 7046 2722 7098
rect 2722 7046 2734 7098
rect 2734 7046 2748 7098
rect 2772 7046 2786 7098
rect 2786 7046 2798 7098
rect 2798 7046 2828 7098
rect 2852 7046 2862 7098
rect 2862 7046 2908 7098
rect 2612 7044 2668 7046
rect 2692 7044 2748 7046
rect 2772 7044 2828 7046
rect 2852 7044 2908 7046
rect 4820 7098 4876 7100
rect 4900 7098 4956 7100
rect 4980 7098 5036 7100
rect 5060 7098 5116 7100
rect 4820 7046 4866 7098
rect 4866 7046 4876 7098
rect 4900 7046 4930 7098
rect 4930 7046 4942 7098
rect 4942 7046 4956 7098
rect 4980 7046 4994 7098
rect 4994 7046 5006 7098
rect 5006 7046 5036 7098
rect 5060 7046 5070 7098
rect 5070 7046 5116 7098
rect 4820 7044 4876 7046
rect 4900 7044 4956 7046
rect 4980 7044 5036 7046
rect 5060 7044 5116 7046
rect 7028 7098 7084 7100
rect 7108 7098 7164 7100
rect 7188 7098 7244 7100
rect 7268 7098 7324 7100
rect 7028 7046 7074 7098
rect 7074 7046 7084 7098
rect 7108 7046 7138 7098
rect 7138 7046 7150 7098
rect 7150 7046 7164 7098
rect 7188 7046 7202 7098
rect 7202 7046 7214 7098
rect 7214 7046 7244 7098
rect 7268 7046 7278 7098
rect 7278 7046 7324 7098
rect 7028 7044 7084 7046
rect 7108 7044 7164 7046
rect 7188 7044 7244 7046
rect 7268 7044 7324 7046
rect 9236 7098 9292 7100
rect 9316 7098 9372 7100
rect 9396 7098 9452 7100
rect 9476 7098 9532 7100
rect 9236 7046 9282 7098
rect 9282 7046 9292 7098
rect 9316 7046 9346 7098
rect 9346 7046 9358 7098
rect 9358 7046 9372 7098
rect 9396 7046 9410 7098
rect 9410 7046 9422 7098
rect 9422 7046 9452 7098
rect 9476 7046 9486 7098
rect 9486 7046 9532 7098
rect 9236 7044 9292 7046
rect 9316 7044 9372 7046
rect 9396 7044 9452 7046
rect 9476 7044 9532 7046
rect 1508 6554 1564 6556
rect 1588 6554 1644 6556
rect 1668 6554 1724 6556
rect 1748 6554 1804 6556
rect 1508 6502 1554 6554
rect 1554 6502 1564 6554
rect 1588 6502 1618 6554
rect 1618 6502 1630 6554
rect 1630 6502 1644 6554
rect 1668 6502 1682 6554
rect 1682 6502 1694 6554
rect 1694 6502 1724 6554
rect 1748 6502 1758 6554
rect 1758 6502 1804 6554
rect 1508 6500 1564 6502
rect 1588 6500 1644 6502
rect 1668 6500 1724 6502
rect 1748 6500 1804 6502
rect 3716 6554 3772 6556
rect 3796 6554 3852 6556
rect 3876 6554 3932 6556
rect 3956 6554 4012 6556
rect 3716 6502 3762 6554
rect 3762 6502 3772 6554
rect 3796 6502 3826 6554
rect 3826 6502 3838 6554
rect 3838 6502 3852 6554
rect 3876 6502 3890 6554
rect 3890 6502 3902 6554
rect 3902 6502 3932 6554
rect 3956 6502 3966 6554
rect 3966 6502 4012 6554
rect 3716 6500 3772 6502
rect 3796 6500 3852 6502
rect 3876 6500 3932 6502
rect 3956 6500 4012 6502
rect 5924 6554 5980 6556
rect 6004 6554 6060 6556
rect 6084 6554 6140 6556
rect 6164 6554 6220 6556
rect 5924 6502 5970 6554
rect 5970 6502 5980 6554
rect 6004 6502 6034 6554
rect 6034 6502 6046 6554
rect 6046 6502 6060 6554
rect 6084 6502 6098 6554
rect 6098 6502 6110 6554
rect 6110 6502 6140 6554
rect 6164 6502 6174 6554
rect 6174 6502 6220 6554
rect 5924 6500 5980 6502
rect 6004 6500 6060 6502
rect 6084 6500 6140 6502
rect 6164 6500 6220 6502
rect 8132 6554 8188 6556
rect 8212 6554 8268 6556
rect 8292 6554 8348 6556
rect 8372 6554 8428 6556
rect 8132 6502 8178 6554
rect 8178 6502 8188 6554
rect 8212 6502 8242 6554
rect 8242 6502 8254 6554
rect 8254 6502 8268 6554
rect 8292 6502 8306 6554
rect 8306 6502 8318 6554
rect 8318 6502 8348 6554
rect 8372 6502 8382 6554
rect 8382 6502 8428 6554
rect 8132 6500 8188 6502
rect 8212 6500 8268 6502
rect 8292 6500 8348 6502
rect 8372 6500 8428 6502
rect 2612 6010 2668 6012
rect 2692 6010 2748 6012
rect 2772 6010 2828 6012
rect 2852 6010 2908 6012
rect 2612 5958 2658 6010
rect 2658 5958 2668 6010
rect 2692 5958 2722 6010
rect 2722 5958 2734 6010
rect 2734 5958 2748 6010
rect 2772 5958 2786 6010
rect 2786 5958 2798 6010
rect 2798 5958 2828 6010
rect 2852 5958 2862 6010
rect 2862 5958 2908 6010
rect 2612 5956 2668 5958
rect 2692 5956 2748 5958
rect 2772 5956 2828 5958
rect 2852 5956 2908 5958
rect 4820 6010 4876 6012
rect 4900 6010 4956 6012
rect 4980 6010 5036 6012
rect 5060 6010 5116 6012
rect 4820 5958 4866 6010
rect 4866 5958 4876 6010
rect 4900 5958 4930 6010
rect 4930 5958 4942 6010
rect 4942 5958 4956 6010
rect 4980 5958 4994 6010
rect 4994 5958 5006 6010
rect 5006 5958 5036 6010
rect 5060 5958 5070 6010
rect 5070 5958 5116 6010
rect 4820 5956 4876 5958
rect 4900 5956 4956 5958
rect 4980 5956 5036 5958
rect 5060 5956 5116 5958
rect 7028 6010 7084 6012
rect 7108 6010 7164 6012
rect 7188 6010 7244 6012
rect 7268 6010 7324 6012
rect 7028 5958 7074 6010
rect 7074 5958 7084 6010
rect 7108 5958 7138 6010
rect 7138 5958 7150 6010
rect 7150 5958 7164 6010
rect 7188 5958 7202 6010
rect 7202 5958 7214 6010
rect 7214 5958 7244 6010
rect 7268 5958 7278 6010
rect 7278 5958 7324 6010
rect 7028 5956 7084 5958
rect 7108 5956 7164 5958
rect 7188 5956 7244 5958
rect 7268 5956 7324 5958
rect 9236 6010 9292 6012
rect 9316 6010 9372 6012
rect 9396 6010 9452 6012
rect 9476 6010 9532 6012
rect 9236 5958 9282 6010
rect 9282 5958 9292 6010
rect 9316 5958 9346 6010
rect 9346 5958 9358 6010
rect 9358 5958 9372 6010
rect 9396 5958 9410 6010
rect 9410 5958 9422 6010
rect 9422 5958 9452 6010
rect 9476 5958 9486 6010
rect 9486 5958 9532 6010
rect 9236 5956 9292 5958
rect 9316 5956 9372 5958
rect 9396 5956 9452 5958
rect 9476 5956 9532 5958
rect 1508 5466 1564 5468
rect 1588 5466 1644 5468
rect 1668 5466 1724 5468
rect 1748 5466 1804 5468
rect 1508 5414 1554 5466
rect 1554 5414 1564 5466
rect 1588 5414 1618 5466
rect 1618 5414 1630 5466
rect 1630 5414 1644 5466
rect 1668 5414 1682 5466
rect 1682 5414 1694 5466
rect 1694 5414 1724 5466
rect 1748 5414 1758 5466
rect 1758 5414 1804 5466
rect 1508 5412 1564 5414
rect 1588 5412 1644 5414
rect 1668 5412 1724 5414
rect 1748 5412 1804 5414
rect 3716 5466 3772 5468
rect 3796 5466 3852 5468
rect 3876 5466 3932 5468
rect 3956 5466 4012 5468
rect 3716 5414 3762 5466
rect 3762 5414 3772 5466
rect 3796 5414 3826 5466
rect 3826 5414 3838 5466
rect 3838 5414 3852 5466
rect 3876 5414 3890 5466
rect 3890 5414 3902 5466
rect 3902 5414 3932 5466
rect 3956 5414 3966 5466
rect 3966 5414 4012 5466
rect 3716 5412 3772 5414
rect 3796 5412 3852 5414
rect 3876 5412 3932 5414
rect 3956 5412 4012 5414
rect 5924 5466 5980 5468
rect 6004 5466 6060 5468
rect 6084 5466 6140 5468
rect 6164 5466 6220 5468
rect 5924 5414 5970 5466
rect 5970 5414 5980 5466
rect 6004 5414 6034 5466
rect 6034 5414 6046 5466
rect 6046 5414 6060 5466
rect 6084 5414 6098 5466
rect 6098 5414 6110 5466
rect 6110 5414 6140 5466
rect 6164 5414 6174 5466
rect 6174 5414 6220 5466
rect 5924 5412 5980 5414
rect 6004 5412 6060 5414
rect 6084 5412 6140 5414
rect 6164 5412 6220 5414
rect 8132 5466 8188 5468
rect 8212 5466 8268 5468
rect 8292 5466 8348 5468
rect 8372 5466 8428 5468
rect 8132 5414 8178 5466
rect 8178 5414 8188 5466
rect 8212 5414 8242 5466
rect 8242 5414 8254 5466
rect 8254 5414 8268 5466
rect 8292 5414 8306 5466
rect 8306 5414 8318 5466
rect 8318 5414 8348 5466
rect 8372 5414 8382 5466
rect 8382 5414 8428 5466
rect 8132 5412 8188 5414
rect 8212 5412 8268 5414
rect 8292 5412 8348 5414
rect 8372 5412 8428 5414
rect 2612 4922 2668 4924
rect 2692 4922 2748 4924
rect 2772 4922 2828 4924
rect 2852 4922 2908 4924
rect 2612 4870 2658 4922
rect 2658 4870 2668 4922
rect 2692 4870 2722 4922
rect 2722 4870 2734 4922
rect 2734 4870 2748 4922
rect 2772 4870 2786 4922
rect 2786 4870 2798 4922
rect 2798 4870 2828 4922
rect 2852 4870 2862 4922
rect 2862 4870 2908 4922
rect 2612 4868 2668 4870
rect 2692 4868 2748 4870
rect 2772 4868 2828 4870
rect 2852 4868 2908 4870
rect 4820 4922 4876 4924
rect 4900 4922 4956 4924
rect 4980 4922 5036 4924
rect 5060 4922 5116 4924
rect 4820 4870 4866 4922
rect 4866 4870 4876 4922
rect 4900 4870 4930 4922
rect 4930 4870 4942 4922
rect 4942 4870 4956 4922
rect 4980 4870 4994 4922
rect 4994 4870 5006 4922
rect 5006 4870 5036 4922
rect 5060 4870 5070 4922
rect 5070 4870 5116 4922
rect 4820 4868 4876 4870
rect 4900 4868 4956 4870
rect 4980 4868 5036 4870
rect 5060 4868 5116 4870
rect 7028 4922 7084 4924
rect 7108 4922 7164 4924
rect 7188 4922 7244 4924
rect 7268 4922 7324 4924
rect 7028 4870 7074 4922
rect 7074 4870 7084 4922
rect 7108 4870 7138 4922
rect 7138 4870 7150 4922
rect 7150 4870 7164 4922
rect 7188 4870 7202 4922
rect 7202 4870 7214 4922
rect 7214 4870 7244 4922
rect 7268 4870 7278 4922
rect 7278 4870 7324 4922
rect 7028 4868 7084 4870
rect 7108 4868 7164 4870
rect 7188 4868 7244 4870
rect 7268 4868 7324 4870
rect 9236 4922 9292 4924
rect 9316 4922 9372 4924
rect 9396 4922 9452 4924
rect 9476 4922 9532 4924
rect 9236 4870 9282 4922
rect 9282 4870 9292 4922
rect 9316 4870 9346 4922
rect 9346 4870 9358 4922
rect 9358 4870 9372 4922
rect 9396 4870 9410 4922
rect 9410 4870 9422 4922
rect 9422 4870 9452 4922
rect 9476 4870 9486 4922
rect 9486 4870 9532 4922
rect 9236 4868 9292 4870
rect 9316 4868 9372 4870
rect 9396 4868 9452 4870
rect 9476 4868 9532 4870
rect 1508 4378 1564 4380
rect 1588 4378 1644 4380
rect 1668 4378 1724 4380
rect 1748 4378 1804 4380
rect 1508 4326 1554 4378
rect 1554 4326 1564 4378
rect 1588 4326 1618 4378
rect 1618 4326 1630 4378
rect 1630 4326 1644 4378
rect 1668 4326 1682 4378
rect 1682 4326 1694 4378
rect 1694 4326 1724 4378
rect 1748 4326 1758 4378
rect 1758 4326 1804 4378
rect 1508 4324 1564 4326
rect 1588 4324 1644 4326
rect 1668 4324 1724 4326
rect 1748 4324 1804 4326
rect 3716 4378 3772 4380
rect 3796 4378 3852 4380
rect 3876 4378 3932 4380
rect 3956 4378 4012 4380
rect 3716 4326 3762 4378
rect 3762 4326 3772 4378
rect 3796 4326 3826 4378
rect 3826 4326 3838 4378
rect 3838 4326 3852 4378
rect 3876 4326 3890 4378
rect 3890 4326 3902 4378
rect 3902 4326 3932 4378
rect 3956 4326 3966 4378
rect 3966 4326 4012 4378
rect 3716 4324 3772 4326
rect 3796 4324 3852 4326
rect 3876 4324 3932 4326
rect 3956 4324 4012 4326
rect 5924 4378 5980 4380
rect 6004 4378 6060 4380
rect 6084 4378 6140 4380
rect 6164 4378 6220 4380
rect 5924 4326 5970 4378
rect 5970 4326 5980 4378
rect 6004 4326 6034 4378
rect 6034 4326 6046 4378
rect 6046 4326 6060 4378
rect 6084 4326 6098 4378
rect 6098 4326 6110 4378
rect 6110 4326 6140 4378
rect 6164 4326 6174 4378
rect 6174 4326 6220 4378
rect 5924 4324 5980 4326
rect 6004 4324 6060 4326
rect 6084 4324 6140 4326
rect 6164 4324 6220 4326
rect 8132 4378 8188 4380
rect 8212 4378 8268 4380
rect 8292 4378 8348 4380
rect 8372 4378 8428 4380
rect 8132 4326 8178 4378
rect 8178 4326 8188 4378
rect 8212 4326 8242 4378
rect 8242 4326 8254 4378
rect 8254 4326 8268 4378
rect 8292 4326 8306 4378
rect 8306 4326 8318 4378
rect 8318 4326 8348 4378
rect 8372 4326 8382 4378
rect 8382 4326 8428 4378
rect 8132 4324 8188 4326
rect 8212 4324 8268 4326
rect 8292 4324 8348 4326
rect 8372 4324 8428 4326
rect 2612 3834 2668 3836
rect 2692 3834 2748 3836
rect 2772 3834 2828 3836
rect 2852 3834 2908 3836
rect 2612 3782 2658 3834
rect 2658 3782 2668 3834
rect 2692 3782 2722 3834
rect 2722 3782 2734 3834
rect 2734 3782 2748 3834
rect 2772 3782 2786 3834
rect 2786 3782 2798 3834
rect 2798 3782 2828 3834
rect 2852 3782 2862 3834
rect 2862 3782 2908 3834
rect 2612 3780 2668 3782
rect 2692 3780 2748 3782
rect 2772 3780 2828 3782
rect 2852 3780 2908 3782
rect 4820 3834 4876 3836
rect 4900 3834 4956 3836
rect 4980 3834 5036 3836
rect 5060 3834 5116 3836
rect 4820 3782 4866 3834
rect 4866 3782 4876 3834
rect 4900 3782 4930 3834
rect 4930 3782 4942 3834
rect 4942 3782 4956 3834
rect 4980 3782 4994 3834
rect 4994 3782 5006 3834
rect 5006 3782 5036 3834
rect 5060 3782 5070 3834
rect 5070 3782 5116 3834
rect 4820 3780 4876 3782
rect 4900 3780 4956 3782
rect 4980 3780 5036 3782
rect 5060 3780 5116 3782
rect 7028 3834 7084 3836
rect 7108 3834 7164 3836
rect 7188 3834 7244 3836
rect 7268 3834 7324 3836
rect 7028 3782 7074 3834
rect 7074 3782 7084 3834
rect 7108 3782 7138 3834
rect 7138 3782 7150 3834
rect 7150 3782 7164 3834
rect 7188 3782 7202 3834
rect 7202 3782 7214 3834
rect 7214 3782 7244 3834
rect 7268 3782 7278 3834
rect 7278 3782 7324 3834
rect 7028 3780 7084 3782
rect 7108 3780 7164 3782
rect 7188 3780 7244 3782
rect 7268 3780 7324 3782
rect 9236 3834 9292 3836
rect 9316 3834 9372 3836
rect 9396 3834 9452 3836
rect 9476 3834 9532 3836
rect 9236 3782 9282 3834
rect 9282 3782 9292 3834
rect 9316 3782 9346 3834
rect 9346 3782 9358 3834
rect 9358 3782 9372 3834
rect 9396 3782 9410 3834
rect 9410 3782 9422 3834
rect 9422 3782 9452 3834
rect 9476 3782 9486 3834
rect 9486 3782 9532 3834
rect 9236 3780 9292 3782
rect 9316 3780 9372 3782
rect 9396 3780 9452 3782
rect 9476 3780 9532 3782
rect 1508 3290 1564 3292
rect 1588 3290 1644 3292
rect 1668 3290 1724 3292
rect 1748 3290 1804 3292
rect 1508 3238 1554 3290
rect 1554 3238 1564 3290
rect 1588 3238 1618 3290
rect 1618 3238 1630 3290
rect 1630 3238 1644 3290
rect 1668 3238 1682 3290
rect 1682 3238 1694 3290
rect 1694 3238 1724 3290
rect 1748 3238 1758 3290
rect 1758 3238 1804 3290
rect 1508 3236 1564 3238
rect 1588 3236 1644 3238
rect 1668 3236 1724 3238
rect 1748 3236 1804 3238
rect 3716 3290 3772 3292
rect 3796 3290 3852 3292
rect 3876 3290 3932 3292
rect 3956 3290 4012 3292
rect 3716 3238 3762 3290
rect 3762 3238 3772 3290
rect 3796 3238 3826 3290
rect 3826 3238 3838 3290
rect 3838 3238 3852 3290
rect 3876 3238 3890 3290
rect 3890 3238 3902 3290
rect 3902 3238 3932 3290
rect 3956 3238 3966 3290
rect 3966 3238 4012 3290
rect 3716 3236 3772 3238
rect 3796 3236 3852 3238
rect 3876 3236 3932 3238
rect 3956 3236 4012 3238
rect 5924 3290 5980 3292
rect 6004 3290 6060 3292
rect 6084 3290 6140 3292
rect 6164 3290 6220 3292
rect 5924 3238 5970 3290
rect 5970 3238 5980 3290
rect 6004 3238 6034 3290
rect 6034 3238 6046 3290
rect 6046 3238 6060 3290
rect 6084 3238 6098 3290
rect 6098 3238 6110 3290
rect 6110 3238 6140 3290
rect 6164 3238 6174 3290
rect 6174 3238 6220 3290
rect 5924 3236 5980 3238
rect 6004 3236 6060 3238
rect 6084 3236 6140 3238
rect 6164 3236 6220 3238
rect 8132 3290 8188 3292
rect 8212 3290 8268 3292
rect 8292 3290 8348 3292
rect 8372 3290 8428 3292
rect 8132 3238 8178 3290
rect 8178 3238 8188 3290
rect 8212 3238 8242 3290
rect 8242 3238 8254 3290
rect 8254 3238 8268 3290
rect 8292 3238 8306 3290
rect 8306 3238 8318 3290
rect 8318 3238 8348 3290
rect 8372 3238 8382 3290
rect 8382 3238 8428 3290
rect 8132 3236 8188 3238
rect 8212 3236 8268 3238
rect 8292 3236 8348 3238
rect 8372 3236 8428 3238
rect 2612 2746 2668 2748
rect 2692 2746 2748 2748
rect 2772 2746 2828 2748
rect 2852 2746 2908 2748
rect 2612 2694 2658 2746
rect 2658 2694 2668 2746
rect 2692 2694 2722 2746
rect 2722 2694 2734 2746
rect 2734 2694 2748 2746
rect 2772 2694 2786 2746
rect 2786 2694 2798 2746
rect 2798 2694 2828 2746
rect 2852 2694 2862 2746
rect 2862 2694 2908 2746
rect 2612 2692 2668 2694
rect 2692 2692 2748 2694
rect 2772 2692 2828 2694
rect 2852 2692 2908 2694
rect 4820 2746 4876 2748
rect 4900 2746 4956 2748
rect 4980 2746 5036 2748
rect 5060 2746 5116 2748
rect 4820 2694 4866 2746
rect 4866 2694 4876 2746
rect 4900 2694 4930 2746
rect 4930 2694 4942 2746
rect 4942 2694 4956 2746
rect 4980 2694 4994 2746
rect 4994 2694 5006 2746
rect 5006 2694 5036 2746
rect 5060 2694 5070 2746
rect 5070 2694 5116 2746
rect 4820 2692 4876 2694
rect 4900 2692 4956 2694
rect 4980 2692 5036 2694
rect 5060 2692 5116 2694
rect 1508 2202 1564 2204
rect 1588 2202 1644 2204
rect 1668 2202 1724 2204
rect 1748 2202 1804 2204
rect 1508 2150 1554 2202
rect 1554 2150 1564 2202
rect 1588 2150 1618 2202
rect 1618 2150 1630 2202
rect 1630 2150 1644 2202
rect 1668 2150 1682 2202
rect 1682 2150 1694 2202
rect 1694 2150 1724 2202
rect 1748 2150 1758 2202
rect 1758 2150 1804 2202
rect 1508 2148 1564 2150
rect 1588 2148 1644 2150
rect 1668 2148 1724 2150
rect 1748 2148 1804 2150
rect 3716 2202 3772 2204
rect 3796 2202 3852 2204
rect 3876 2202 3932 2204
rect 3956 2202 4012 2204
rect 3716 2150 3762 2202
rect 3762 2150 3772 2202
rect 3796 2150 3826 2202
rect 3826 2150 3838 2202
rect 3838 2150 3852 2202
rect 3876 2150 3890 2202
rect 3890 2150 3902 2202
rect 3902 2150 3932 2202
rect 3956 2150 3966 2202
rect 3966 2150 4012 2202
rect 3716 2148 3772 2150
rect 3796 2148 3852 2150
rect 3876 2148 3932 2150
rect 3956 2148 4012 2150
rect 2612 1658 2668 1660
rect 2692 1658 2748 1660
rect 2772 1658 2828 1660
rect 2852 1658 2908 1660
rect 2612 1606 2658 1658
rect 2658 1606 2668 1658
rect 2692 1606 2722 1658
rect 2722 1606 2734 1658
rect 2734 1606 2748 1658
rect 2772 1606 2786 1658
rect 2786 1606 2798 1658
rect 2798 1606 2828 1658
rect 2852 1606 2862 1658
rect 2862 1606 2908 1658
rect 2612 1604 2668 1606
rect 2692 1604 2748 1606
rect 2772 1604 2828 1606
rect 2852 1604 2908 1606
rect 1508 1114 1564 1116
rect 1588 1114 1644 1116
rect 1668 1114 1724 1116
rect 1748 1114 1804 1116
rect 1508 1062 1554 1114
rect 1554 1062 1564 1114
rect 1588 1062 1618 1114
rect 1618 1062 1630 1114
rect 1630 1062 1644 1114
rect 1668 1062 1682 1114
rect 1682 1062 1694 1114
rect 1694 1062 1724 1114
rect 1748 1062 1758 1114
rect 1758 1062 1804 1114
rect 1508 1060 1564 1062
rect 1588 1060 1644 1062
rect 1668 1060 1724 1062
rect 1748 1060 1804 1062
rect 3716 1114 3772 1116
rect 3796 1114 3852 1116
rect 3876 1114 3932 1116
rect 3956 1114 4012 1116
rect 3716 1062 3762 1114
rect 3762 1062 3772 1114
rect 3796 1062 3826 1114
rect 3826 1062 3838 1114
rect 3838 1062 3852 1114
rect 3876 1062 3890 1114
rect 3890 1062 3902 1114
rect 3902 1062 3932 1114
rect 3956 1062 3966 1114
rect 3966 1062 4012 1114
rect 3716 1060 3772 1062
rect 3796 1060 3852 1062
rect 3876 1060 3932 1062
rect 3956 1060 4012 1062
rect 4820 1658 4876 1660
rect 4900 1658 4956 1660
rect 4980 1658 5036 1660
rect 5060 1658 5116 1660
rect 4820 1606 4866 1658
rect 4866 1606 4876 1658
rect 4900 1606 4930 1658
rect 4930 1606 4942 1658
rect 4942 1606 4956 1658
rect 4980 1606 4994 1658
rect 4994 1606 5006 1658
rect 5006 1606 5036 1658
rect 5060 1606 5070 1658
rect 5070 1606 5116 1658
rect 4820 1604 4876 1606
rect 4900 1604 4956 1606
rect 4980 1604 5036 1606
rect 5060 1604 5116 1606
rect 7028 2746 7084 2748
rect 7108 2746 7164 2748
rect 7188 2746 7244 2748
rect 7268 2746 7324 2748
rect 7028 2694 7074 2746
rect 7074 2694 7084 2746
rect 7108 2694 7138 2746
rect 7138 2694 7150 2746
rect 7150 2694 7164 2746
rect 7188 2694 7202 2746
rect 7202 2694 7214 2746
rect 7214 2694 7244 2746
rect 7268 2694 7278 2746
rect 7278 2694 7324 2746
rect 7028 2692 7084 2694
rect 7108 2692 7164 2694
rect 7188 2692 7244 2694
rect 7268 2692 7324 2694
rect 9236 2746 9292 2748
rect 9316 2746 9372 2748
rect 9396 2746 9452 2748
rect 9476 2746 9532 2748
rect 9236 2694 9282 2746
rect 9282 2694 9292 2746
rect 9316 2694 9346 2746
rect 9346 2694 9358 2746
rect 9358 2694 9372 2746
rect 9396 2694 9410 2746
rect 9410 2694 9422 2746
rect 9422 2694 9452 2746
rect 9476 2694 9486 2746
rect 9486 2694 9532 2746
rect 9236 2692 9292 2694
rect 9316 2692 9372 2694
rect 9396 2692 9452 2694
rect 9476 2692 9532 2694
rect 5924 2202 5980 2204
rect 6004 2202 6060 2204
rect 6084 2202 6140 2204
rect 6164 2202 6220 2204
rect 5924 2150 5970 2202
rect 5970 2150 5980 2202
rect 6004 2150 6034 2202
rect 6034 2150 6046 2202
rect 6046 2150 6060 2202
rect 6084 2150 6098 2202
rect 6098 2150 6110 2202
rect 6110 2150 6140 2202
rect 6164 2150 6174 2202
rect 6174 2150 6220 2202
rect 5924 2148 5980 2150
rect 6004 2148 6060 2150
rect 6084 2148 6140 2150
rect 6164 2148 6220 2150
rect 2612 570 2668 572
rect 2692 570 2748 572
rect 2772 570 2828 572
rect 2852 570 2908 572
rect 2612 518 2658 570
rect 2658 518 2668 570
rect 2692 518 2722 570
rect 2722 518 2734 570
rect 2734 518 2748 570
rect 2772 518 2786 570
rect 2786 518 2798 570
rect 2798 518 2828 570
rect 2852 518 2862 570
rect 2862 518 2908 570
rect 2612 516 2668 518
rect 2692 516 2748 518
rect 2772 516 2828 518
rect 2852 516 2908 518
rect 4820 570 4876 572
rect 4900 570 4956 572
rect 4980 570 5036 572
rect 5060 570 5116 572
rect 4820 518 4866 570
rect 4866 518 4876 570
rect 4900 518 4930 570
rect 4930 518 4942 570
rect 4942 518 4956 570
rect 4980 518 4994 570
rect 4994 518 5006 570
rect 5006 518 5036 570
rect 5060 518 5070 570
rect 5070 518 5116 570
rect 4820 516 4876 518
rect 4900 516 4956 518
rect 4980 516 5036 518
rect 5060 516 5116 518
rect 5924 1114 5980 1116
rect 6004 1114 6060 1116
rect 6084 1114 6140 1116
rect 6164 1114 6220 1116
rect 5924 1062 5970 1114
rect 5970 1062 5980 1114
rect 6004 1062 6034 1114
rect 6034 1062 6046 1114
rect 6046 1062 6060 1114
rect 6084 1062 6098 1114
rect 6098 1062 6110 1114
rect 6110 1062 6140 1114
rect 6164 1062 6174 1114
rect 6174 1062 6220 1114
rect 5924 1060 5980 1062
rect 6004 1060 6060 1062
rect 6084 1060 6140 1062
rect 6164 1060 6220 1062
rect 7028 1658 7084 1660
rect 7108 1658 7164 1660
rect 7188 1658 7244 1660
rect 7268 1658 7324 1660
rect 7028 1606 7074 1658
rect 7074 1606 7084 1658
rect 7108 1606 7138 1658
rect 7138 1606 7150 1658
rect 7150 1606 7164 1658
rect 7188 1606 7202 1658
rect 7202 1606 7214 1658
rect 7214 1606 7244 1658
rect 7268 1606 7278 1658
rect 7278 1606 7324 1658
rect 7028 1604 7084 1606
rect 7108 1604 7164 1606
rect 7188 1604 7244 1606
rect 7268 1604 7324 1606
rect 7028 570 7084 572
rect 7108 570 7164 572
rect 7188 570 7244 572
rect 7268 570 7324 572
rect 7028 518 7074 570
rect 7074 518 7084 570
rect 7108 518 7138 570
rect 7138 518 7150 570
rect 7150 518 7164 570
rect 7188 518 7202 570
rect 7202 518 7214 570
rect 7214 518 7244 570
rect 7268 518 7278 570
rect 7278 518 7324 570
rect 7028 516 7084 518
rect 7108 516 7164 518
rect 7188 516 7244 518
rect 7268 516 7324 518
rect 8132 2202 8188 2204
rect 8212 2202 8268 2204
rect 8292 2202 8348 2204
rect 8372 2202 8428 2204
rect 8132 2150 8178 2202
rect 8178 2150 8188 2202
rect 8212 2150 8242 2202
rect 8242 2150 8254 2202
rect 8254 2150 8268 2202
rect 8292 2150 8306 2202
rect 8306 2150 8318 2202
rect 8318 2150 8348 2202
rect 8372 2150 8382 2202
rect 8382 2150 8428 2202
rect 8132 2148 8188 2150
rect 8212 2148 8268 2150
rect 8292 2148 8348 2150
rect 8372 2148 8428 2150
rect 8132 1114 8188 1116
rect 8212 1114 8268 1116
rect 8292 1114 8348 1116
rect 8372 1114 8428 1116
rect 8132 1062 8178 1114
rect 8178 1062 8188 1114
rect 8212 1062 8242 1114
rect 8242 1062 8254 1114
rect 8254 1062 8268 1114
rect 8292 1062 8306 1114
rect 8306 1062 8318 1114
rect 8318 1062 8348 1114
rect 8372 1062 8382 1114
rect 8382 1062 8428 1114
rect 8132 1060 8188 1062
rect 8212 1060 8268 1062
rect 8292 1060 8348 1062
rect 8372 1060 8428 1062
rect 9236 1658 9292 1660
rect 9316 1658 9372 1660
rect 9396 1658 9452 1660
rect 9476 1658 9532 1660
rect 9236 1606 9282 1658
rect 9282 1606 9292 1658
rect 9316 1606 9346 1658
rect 9346 1606 9358 1658
rect 9358 1606 9372 1658
rect 9396 1606 9410 1658
rect 9410 1606 9422 1658
rect 9422 1606 9452 1658
rect 9476 1606 9486 1658
rect 9486 1606 9532 1658
rect 9236 1604 9292 1606
rect 9316 1604 9372 1606
rect 9396 1604 9452 1606
rect 9476 1604 9532 1606
rect 9236 570 9292 572
rect 9316 570 9372 572
rect 9396 570 9452 572
rect 9476 570 9532 572
rect 9236 518 9282 570
rect 9282 518 9292 570
rect 9316 518 9346 570
rect 9346 518 9358 570
rect 9358 518 9372 570
rect 9396 518 9410 570
rect 9410 518 9422 570
rect 9422 518 9452 570
rect 9476 518 9486 570
rect 9486 518 9532 570
rect 9236 516 9292 518
rect 9316 516 9372 518
rect 9396 516 9452 518
rect 9476 516 9532 518
<< metal3 >>
rect 2602 9280 2918 9281
rect 2602 9216 2608 9280
rect 2672 9216 2688 9280
rect 2752 9216 2768 9280
rect 2832 9216 2848 9280
rect 2912 9216 2918 9280
rect 2602 9215 2918 9216
rect 4810 9280 5126 9281
rect 4810 9216 4816 9280
rect 4880 9216 4896 9280
rect 4960 9216 4976 9280
rect 5040 9216 5056 9280
rect 5120 9216 5126 9280
rect 4810 9215 5126 9216
rect 7018 9280 7334 9281
rect 7018 9216 7024 9280
rect 7088 9216 7104 9280
rect 7168 9216 7184 9280
rect 7248 9216 7264 9280
rect 7328 9216 7334 9280
rect 7018 9215 7334 9216
rect 9226 9280 9542 9281
rect 9226 9216 9232 9280
rect 9296 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9542 9280
rect 9226 9215 9542 9216
rect 1498 8736 1814 8737
rect 1498 8672 1504 8736
rect 1568 8672 1584 8736
rect 1648 8672 1664 8736
rect 1728 8672 1744 8736
rect 1808 8672 1814 8736
rect 1498 8671 1814 8672
rect 3706 8736 4022 8737
rect 3706 8672 3712 8736
rect 3776 8672 3792 8736
rect 3856 8672 3872 8736
rect 3936 8672 3952 8736
rect 4016 8672 4022 8736
rect 3706 8671 4022 8672
rect 5914 8736 6230 8737
rect 5914 8672 5920 8736
rect 5984 8672 6000 8736
rect 6064 8672 6080 8736
rect 6144 8672 6160 8736
rect 6224 8672 6230 8736
rect 5914 8671 6230 8672
rect 8122 8736 8438 8737
rect 8122 8672 8128 8736
rect 8192 8672 8208 8736
rect 8272 8672 8288 8736
rect 8352 8672 8368 8736
rect 8432 8672 8438 8736
rect 8122 8671 8438 8672
rect 2602 8192 2918 8193
rect 2602 8128 2608 8192
rect 2672 8128 2688 8192
rect 2752 8128 2768 8192
rect 2832 8128 2848 8192
rect 2912 8128 2918 8192
rect 2602 8127 2918 8128
rect 4810 8192 5126 8193
rect 4810 8128 4816 8192
rect 4880 8128 4896 8192
rect 4960 8128 4976 8192
rect 5040 8128 5056 8192
rect 5120 8128 5126 8192
rect 4810 8127 5126 8128
rect 7018 8192 7334 8193
rect 7018 8128 7024 8192
rect 7088 8128 7104 8192
rect 7168 8128 7184 8192
rect 7248 8128 7264 8192
rect 7328 8128 7334 8192
rect 7018 8127 7334 8128
rect 9226 8192 9542 8193
rect 9226 8128 9232 8192
rect 9296 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9542 8192
rect 9226 8127 9542 8128
rect 1498 7648 1814 7649
rect 1498 7584 1504 7648
rect 1568 7584 1584 7648
rect 1648 7584 1664 7648
rect 1728 7584 1744 7648
rect 1808 7584 1814 7648
rect 1498 7583 1814 7584
rect 3706 7648 4022 7649
rect 3706 7584 3712 7648
rect 3776 7584 3792 7648
rect 3856 7584 3872 7648
rect 3936 7584 3952 7648
rect 4016 7584 4022 7648
rect 3706 7583 4022 7584
rect 5914 7648 6230 7649
rect 5914 7584 5920 7648
rect 5984 7584 6000 7648
rect 6064 7584 6080 7648
rect 6144 7584 6160 7648
rect 6224 7584 6230 7648
rect 5914 7583 6230 7584
rect 8122 7648 8438 7649
rect 8122 7584 8128 7648
rect 8192 7584 8208 7648
rect 8272 7584 8288 7648
rect 8352 7584 8368 7648
rect 8432 7584 8438 7648
rect 8122 7583 8438 7584
rect 2602 7104 2918 7105
rect 2602 7040 2608 7104
rect 2672 7040 2688 7104
rect 2752 7040 2768 7104
rect 2832 7040 2848 7104
rect 2912 7040 2918 7104
rect 2602 7039 2918 7040
rect 4810 7104 5126 7105
rect 4810 7040 4816 7104
rect 4880 7040 4896 7104
rect 4960 7040 4976 7104
rect 5040 7040 5056 7104
rect 5120 7040 5126 7104
rect 4810 7039 5126 7040
rect 7018 7104 7334 7105
rect 7018 7040 7024 7104
rect 7088 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7334 7104
rect 7018 7039 7334 7040
rect 9226 7104 9542 7105
rect 9226 7040 9232 7104
rect 9296 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9542 7104
rect 9226 7039 9542 7040
rect 1498 6560 1814 6561
rect 1498 6496 1504 6560
rect 1568 6496 1584 6560
rect 1648 6496 1664 6560
rect 1728 6496 1744 6560
rect 1808 6496 1814 6560
rect 1498 6495 1814 6496
rect 3706 6560 4022 6561
rect 3706 6496 3712 6560
rect 3776 6496 3792 6560
rect 3856 6496 3872 6560
rect 3936 6496 3952 6560
rect 4016 6496 4022 6560
rect 3706 6495 4022 6496
rect 5914 6560 6230 6561
rect 5914 6496 5920 6560
rect 5984 6496 6000 6560
rect 6064 6496 6080 6560
rect 6144 6496 6160 6560
rect 6224 6496 6230 6560
rect 5914 6495 6230 6496
rect 8122 6560 8438 6561
rect 8122 6496 8128 6560
rect 8192 6496 8208 6560
rect 8272 6496 8288 6560
rect 8352 6496 8368 6560
rect 8432 6496 8438 6560
rect 8122 6495 8438 6496
rect 2602 6016 2918 6017
rect 2602 5952 2608 6016
rect 2672 5952 2688 6016
rect 2752 5952 2768 6016
rect 2832 5952 2848 6016
rect 2912 5952 2918 6016
rect 2602 5951 2918 5952
rect 4810 6016 5126 6017
rect 4810 5952 4816 6016
rect 4880 5952 4896 6016
rect 4960 5952 4976 6016
rect 5040 5952 5056 6016
rect 5120 5952 5126 6016
rect 4810 5951 5126 5952
rect 7018 6016 7334 6017
rect 7018 5952 7024 6016
rect 7088 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7334 6016
rect 7018 5951 7334 5952
rect 9226 6016 9542 6017
rect 9226 5952 9232 6016
rect 9296 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9542 6016
rect 9226 5951 9542 5952
rect 1498 5472 1814 5473
rect 1498 5408 1504 5472
rect 1568 5408 1584 5472
rect 1648 5408 1664 5472
rect 1728 5408 1744 5472
rect 1808 5408 1814 5472
rect 1498 5407 1814 5408
rect 3706 5472 4022 5473
rect 3706 5408 3712 5472
rect 3776 5408 3792 5472
rect 3856 5408 3872 5472
rect 3936 5408 3952 5472
rect 4016 5408 4022 5472
rect 3706 5407 4022 5408
rect 5914 5472 6230 5473
rect 5914 5408 5920 5472
rect 5984 5408 6000 5472
rect 6064 5408 6080 5472
rect 6144 5408 6160 5472
rect 6224 5408 6230 5472
rect 5914 5407 6230 5408
rect 8122 5472 8438 5473
rect 8122 5408 8128 5472
rect 8192 5408 8208 5472
rect 8272 5408 8288 5472
rect 8352 5408 8368 5472
rect 8432 5408 8438 5472
rect 8122 5407 8438 5408
rect 2602 4928 2918 4929
rect 2602 4864 2608 4928
rect 2672 4864 2688 4928
rect 2752 4864 2768 4928
rect 2832 4864 2848 4928
rect 2912 4864 2918 4928
rect 2602 4863 2918 4864
rect 4810 4928 5126 4929
rect 4810 4864 4816 4928
rect 4880 4864 4896 4928
rect 4960 4864 4976 4928
rect 5040 4864 5056 4928
rect 5120 4864 5126 4928
rect 4810 4863 5126 4864
rect 7018 4928 7334 4929
rect 7018 4864 7024 4928
rect 7088 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7334 4928
rect 7018 4863 7334 4864
rect 9226 4928 9542 4929
rect 9226 4864 9232 4928
rect 9296 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9542 4928
rect 9226 4863 9542 4864
rect 1498 4384 1814 4385
rect 1498 4320 1504 4384
rect 1568 4320 1584 4384
rect 1648 4320 1664 4384
rect 1728 4320 1744 4384
rect 1808 4320 1814 4384
rect 1498 4319 1814 4320
rect 3706 4384 4022 4385
rect 3706 4320 3712 4384
rect 3776 4320 3792 4384
rect 3856 4320 3872 4384
rect 3936 4320 3952 4384
rect 4016 4320 4022 4384
rect 3706 4319 4022 4320
rect 5914 4384 6230 4385
rect 5914 4320 5920 4384
rect 5984 4320 6000 4384
rect 6064 4320 6080 4384
rect 6144 4320 6160 4384
rect 6224 4320 6230 4384
rect 5914 4319 6230 4320
rect 8122 4384 8438 4385
rect 8122 4320 8128 4384
rect 8192 4320 8208 4384
rect 8272 4320 8288 4384
rect 8352 4320 8368 4384
rect 8432 4320 8438 4384
rect 8122 4319 8438 4320
rect 2602 3840 2918 3841
rect 2602 3776 2608 3840
rect 2672 3776 2688 3840
rect 2752 3776 2768 3840
rect 2832 3776 2848 3840
rect 2912 3776 2918 3840
rect 2602 3775 2918 3776
rect 4810 3840 5126 3841
rect 4810 3776 4816 3840
rect 4880 3776 4896 3840
rect 4960 3776 4976 3840
rect 5040 3776 5056 3840
rect 5120 3776 5126 3840
rect 4810 3775 5126 3776
rect 7018 3840 7334 3841
rect 7018 3776 7024 3840
rect 7088 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7334 3840
rect 7018 3775 7334 3776
rect 9226 3840 9542 3841
rect 9226 3776 9232 3840
rect 9296 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9542 3840
rect 9226 3775 9542 3776
rect 1498 3296 1814 3297
rect 1498 3232 1504 3296
rect 1568 3232 1584 3296
rect 1648 3232 1664 3296
rect 1728 3232 1744 3296
rect 1808 3232 1814 3296
rect 1498 3231 1814 3232
rect 3706 3296 4022 3297
rect 3706 3232 3712 3296
rect 3776 3232 3792 3296
rect 3856 3232 3872 3296
rect 3936 3232 3952 3296
rect 4016 3232 4022 3296
rect 3706 3231 4022 3232
rect 5914 3296 6230 3297
rect 5914 3232 5920 3296
rect 5984 3232 6000 3296
rect 6064 3232 6080 3296
rect 6144 3232 6160 3296
rect 6224 3232 6230 3296
rect 5914 3231 6230 3232
rect 8122 3296 8438 3297
rect 8122 3232 8128 3296
rect 8192 3232 8208 3296
rect 8272 3232 8288 3296
rect 8352 3232 8368 3296
rect 8432 3232 8438 3296
rect 8122 3231 8438 3232
rect 2602 2752 2918 2753
rect 2602 2688 2608 2752
rect 2672 2688 2688 2752
rect 2752 2688 2768 2752
rect 2832 2688 2848 2752
rect 2912 2688 2918 2752
rect 2602 2687 2918 2688
rect 4810 2752 5126 2753
rect 4810 2688 4816 2752
rect 4880 2688 4896 2752
rect 4960 2688 4976 2752
rect 5040 2688 5056 2752
rect 5120 2688 5126 2752
rect 4810 2687 5126 2688
rect 7018 2752 7334 2753
rect 7018 2688 7024 2752
rect 7088 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7334 2752
rect 7018 2687 7334 2688
rect 9226 2752 9542 2753
rect 9226 2688 9232 2752
rect 9296 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9542 2752
rect 9226 2687 9542 2688
rect 1498 2208 1814 2209
rect 1498 2144 1504 2208
rect 1568 2144 1584 2208
rect 1648 2144 1664 2208
rect 1728 2144 1744 2208
rect 1808 2144 1814 2208
rect 1498 2143 1814 2144
rect 3706 2208 4022 2209
rect 3706 2144 3712 2208
rect 3776 2144 3792 2208
rect 3856 2144 3872 2208
rect 3936 2144 3952 2208
rect 4016 2144 4022 2208
rect 3706 2143 4022 2144
rect 5914 2208 6230 2209
rect 5914 2144 5920 2208
rect 5984 2144 6000 2208
rect 6064 2144 6080 2208
rect 6144 2144 6160 2208
rect 6224 2144 6230 2208
rect 5914 2143 6230 2144
rect 8122 2208 8438 2209
rect 8122 2144 8128 2208
rect 8192 2144 8208 2208
rect 8272 2144 8288 2208
rect 8352 2144 8368 2208
rect 8432 2144 8438 2208
rect 8122 2143 8438 2144
rect 2602 1664 2918 1665
rect 2602 1600 2608 1664
rect 2672 1600 2688 1664
rect 2752 1600 2768 1664
rect 2832 1600 2848 1664
rect 2912 1600 2918 1664
rect 2602 1599 2918 1600
rect 4810 1664 5126 1665
rect 4810 1600 4816 1664
rect 4880 1600 4896 1664
rect 4960 1600 4976 1664
rect 5040 1600 5056 1664
rect 5120 1600 5126 1664
rect 4810 1599 5126 1600
rect 7018 1664 7334 1665
rect 7018 1600 7024 1664
rect 7088 1600 7104 1664
rect 7168 1600 7184 1664
rect 7248 1600 7264 1664
rect 7328 1600 7334 1664
rect 7018 1599 7334 1600
rect 9226 1664 9542 1665
rect 9226 1600 9232 1664
rect 9296 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9542 1664
rect 9226 1599 9542 1600
rect 1498 1120 1814 1121
rect 1498 1056 1504 1120
rect 1568 1056 1584 1120
rect 1648 1056 1664 1120
rect 1728 1056 1744 1120
rect 1808 1056 1814 1120
rect 1498 1055 1814 1056
rect 3706 1120 4022 1121
rect 3706 1056 3712 1120
rect 3776 1056 3792 1120
rect 3856 1056 3872 1120
rect 3936 1056 3952 1120
rect 4016 1056 4022 1120
rect 3706 1055 4022 1056
rect 5914 1120 6230 1121
rect 5914 1056 5920 1120
rect 5984 1056 6000 1120
rect 6064 1056 6080 1120
rect 6144 1056 6160 1120
rect 6224 1056 6230 1120
rect 5914 1055 6230 1056
rect 8122 1120 8438 1121
rect 8122 1056 8128 1120
rect 8192 1056 8208 1120
rect 8272 1056 8288 1120
rect 8352 1056 8368 1120
rect 8432 1056 8438 1120
rect 8122 1055 8438 1056
rect 2602 576 2918 577
rect 2602 512 2608 576
rect 2672 512 2688 576
rect 2752 512 2768 576
rect 2832 512 2848 576
rect 2912 512 2918 576
rect 2602 511 2918 512
rect 4810 576 5126 577
rect 4810 512 4816 576
rect 4880 512 4896 576
rect 4960 512 4976 576
rect 5040 512 5056 576
rect 5120 512 5126 576
rect 4810 511 5126 512
rect 7018 576 7334 577
rect 7018 512 7024 576
rect 7088 512 7104 576
rect 7168 512 7184 576
rect 7248 512 7264 576
rect 7328 512 7334 576
rect 7018 511 7334 512
rect 9226 576 9542 577
rect 9226 512 9232 576
rect 9296 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9542 576
rect 9226 511 9542 512
<< via3 >>
rect 2608 9276 2672 9280
rect 2608 9220 2612 9276
rect 2612 9220 2668 9276
rect 2668 9220 2672 9276
rect 2608 9216 2672 9220
rect 2688 9276 2752 9280
rect 2688 9220 2692 9276
rect 2692 9220 2748 9276
rect 2748 9220 2752 9276
rect 2688 9216 2752 9220
rect 2768 9276 2832 9280
rect 2768 9220 2772 9276
rect 2772 9220 2828 9276
rect 2828 9220 2832 9276
rect 2768 9216 2832 9220
rect 2848 9276 2912 9280
rect 2848 9220 2852 9276
rect 2852 9220 2908 9276
rect 2908 9220 2912 9276
rect 2848 9216 2912 9220
rect 4816 9276 4880 9280
rect 4816 9220 4820 9276
rect 4820 9220 4876 9276
rect 4876 9220 4880 9276
rect 4816 9216 4880 9220
rect 4896 9276 4960 9280
rect 4896 9220 4900 9276
rect 4900 9220 4956 9276
rect 4956 9220 4960 9276
rect 4896 9216 4960 9220
rect 4976 9276 5040 9280
rect 4976 9220 4980 9276
rect 4980 9220 5036 9276
rect 5036 9220 5040 9276
rect 4976 9216 5040 9220
rect 5056 9276 5120 9280
rect 5056 9220 5060 9276
rect 5060 9220 5116 9276
rect 5116 9220 5120 9276
rect 5056 9216 5120 9220
rect 7024 9276 7088 9280
rect 7024 9220 7028 9276
rect 7028 9220 7084 9276
rect 7084 9220 7088 9276
rect 7024 9216 7088 9220
rect 7104 9276 7168 9280
rect 7104 9220 7108 9276
rect 7108 9220 7164 9276
rect 7164 9220 7168 9276
rect 7104 9216 7168 9220
rect 7184 9276 7248 9280
rect 7184 9220 7188 9276
rect 7188 9220 7244 9276
rect 7244 9220 7248 9276
rect 7184 9216 7248 9220
rect 7264 9276 7328 9280
rect 7264 9220 7268 9276
rect 7268 9220 7324 9276
rect 7324 9220 7328 9276
rect 7264 9216 7328 9220
rect 9232 9276 9296 9280
rect 9232 9220 9236 9276
rect 9236 9220 9292 9276
rect 9292 9220 9296 9276
rect 9232 9216 9296 9220
rect 9312 9276 9376 9280
rect 9312 9220 9316 9276
rect 9316 9220 9372 9276
rect 9372 9220 9376 9276
rect 9312 9216 9376 9220
rect 9392 9276 9456 9280
rect 9392 9220 9396 9276
rect 9396 9220 9452 9276
rect 9452 9220 9456 9276
rect 9392 9216 9456 9220
rect 9472 9276 9536 9280
rect 9472 9220 9476 9276
rect 9476 9220 9532 9276
rect 9532 9220 9536 9276
rect 9472 9216 9536 9220
rect 1504 8732 1568 8736
rect 1504 8676 1508 8732
rect 1508 8676 1564 8732
rect 1564 8676 1568 8732
rect 1504 8672 1568 8676
rect 1584 8732 1648 8736
rect 1584 8676 1588 8732
rect 1588 8676 1644 8732
rect 1644 8676 1648 8732
rect 1584 8672 1648 8676
rect 1664 8732 1728 8736
rect 1664 8676 1668 8732
rect 1668 8676 1724 8732
rect 1724 8676 1728 8732
rect 1664 8672 1728 8676
rect 1744 8732 1808 8736
rect 1744 8676 1748 8732
rect 1748 8676 1804 8732
rect 1804 8676 1808 8732
rect 1744 8672 1808 8676
rect 3712 8732 3776 8736
rect 3712 8676 3716 8732
rect 3716 8676 3772 8732
rect 3772 8676 3776 8732
rect 3712 8672 3776 8676
rect 3792 8732 3856 8736
rect 3792 8676 3796 8732
rect 3796 8676 3852 8732
rect 3852 8676 3856 8732
rect 3792 8672 3856 8676
rect 3872 8732 3936 8736
rect 3872 8676 3876 8732
rect 3876 8676 3932 8732
rect 3932 8676 3936 8732
rect 3872 8672 3936 8676
rect 3952 8732 4016 8736
rect 3952 8676 3956 8732
rect 3956 8676 4012 8732
rect 4012 8676 4016 8732
rect 3952 8672 4016 8676
rect 5920 8732 5984 8736
rect 5920 8676 5924 8732
rect 5924 8676 5980 8732
rect 5980 8676 5984 8732
rect 5920 8672 5984 8676
rect 6000 8732 6064 8736
rect 6000 8676 6004 8732
rect 6004 8676 6060 8732
rect 6060 8676 6064 8732
rect 6000 8672 6064 8676
rect 6080 8732 6144 8736
rect 6080 8676 6084 8732
rect 6084 8676 6140 8732
rect 6140 8676 6144 8732
rect 6080 8672 6144 8676
rect 6160 8732 6224 8736
rect 6160 8676 6164 8732
rect 6164 8676 6220 8732
rect 6220 8676 6224 8732
rect 6160 8672 6224 8676
rect 8128 8732 8192 8736
rect 8128 8676 8132 8732
rect 8132 8676 8188 8732
rect 8188 8676 8192 8732
rect 8128 8672 8192 8676
rect 8208 8732 8272 8736
rect 8208 8676 8212 8732
rect 8212 8676 8268 8732
rect 8268 8676 8272 8732
rect 8208 8672 8272 8676
rect 8288 8732 8352 8736
rect 8288 8676 8292 8732
rect 8292 8676 8348 8732
rect 8348 8676 8352 8732
rect 8288 8672 8352 8676
rect 8368 8732 8432 8736
rect 8368 8676 8372 8732
rect 8372 8676 8428 8732
rect 8428 8676 8432 8732
rect 8368 8672 8432 8676
rect 2608 8188 2672 8192
rect 2608 8132 2612 8188
rect 2612 8132 2668 8188
rect 2668 8132 2672 8188
rect 2608 8128 2672 8132
rect 2688 8188 2752 8192
rect 2688 8132 2692 8188
rect 2692 8132 2748 8188
rect 2748 8132 2752 8188
rect 2688 8128 2752 8132
rect 2768 8188 2832 8192
rect 2768 8132 2772 8188
rect 2772 8132 2828 8188
rect 2828 8132 2832 8188
rect 2768 8128 2832 8132
rect 2848 8188 2912 8192
rect 2848 8132 2852 8188
rect 2852 8132 2908 8188
rect 2908 8132 2912 8188
rect 2848 8128 2912 8132
rect 4816 8188 4880 8192
rect 4816 8132 4820 8188
rect 4820 8132 4876 8188
rect 4876 8132 4880 8188
rect 4816 8128 4880 8132
rect 4896 8188 4960 8192
rect 4896 8132 4900 8188
rect 4900 8132 4956 8188
rect 4956 8132 4960 8188
rect 4896 8128 4960 8132
rect 4976 8188 5040 8192
rect 4976 8132 4980 8188
rect 4980 8132 5036 8188
rect 5036 8132 5040 8188
rect 4976 8128 5040 8132
rect 5056 8188 5120 8192
rect 5056 8132 5060 8188
rect 5060 8132 5116 8188
rect 5116 8132 5120 8188
rect 5056 8128 5120 8132
rect 7024 8188 7088 8192
rect 7024 8132 7028 8188
rect 7028 8132 7084 8188
rect 7084 8132 7088 8188
rect 7024 8128 7088 8132
rect 7104 8188 7168 8192
rect 7104 8132 7108 8188
rect 7108 8132 7164 8188
rect 7164 8132 7168 8188
rect 7104 8128 7168 8132
rect 7184 8188 7248 8192
rect 7184 8132 7188 8188
rect 7188 8132 7244 8188
rect 7244 8132 7248 8188
rect 7184 8128 7248 8132
rect 7264 8188 7328 8192
rect 7264 8132 7268 8188
rect 7268 8132 7324 8188
rect 7324 8132 7328 8188
rect 7264 8128 7328 8132
rect 9232 8188 9296 8192
rect 9232 8132 9236 8188
rect 9236 8132 9292 8188
rect 9292 8132 9296 8188
rect 9232 8128 9296 8132
rect 9312 8188 9376 8192
rect 9312 8132 9316 8188
rect 9316 8132 9372 8188
rect 9372 8132 9376 8188
rect 9312 8128 9376 8132
rect 9392 8188 9456 8192
rect 9392 8132 9396 8188
rect 9396 8132 9452 8188
rect 9452 8132 9456 8188
rect 9392 8128 9456 8132
rect 9472 8188 9536 8192
rect 9472 8132 9476 8188
rect 9476 8132 9532 8188
rect 9532 8132 9536 8188
rect 9472 8128 9536 8132
rect 1504 7644 1568 7648
rect 1504 7588 1508 7644
rect 1508 7588 1564 7644
rect 1564 7588 1568 7644
rect 1504 7584 1568 7588
rect 1584 7644 1648 7648
rect 1584 7588 1588 7644
rect 1588 7588 1644 7644
rect 1644 7588 1648 7644
rect 1584 7584 1648 7588
rect 1664 7644 1728 7648
rect 1664 7588 1668 7644
rect 1668 7588 1724 7644
rect 1724 7588 1728 7644
rect 1664 7584 1728 7588
rect 1744 7644 1808 7648
rect 1744 7588 1748 7644
rect 1748 7588 1804 7644
rect 1804 7588 1808 7644
rect 1744 7584 1808 7588
rect 3712 7644 3776 7648
rect 3712 7588 3716 7644
rect 3716 7588 3772 7644
rect 3772 7588 3776 7644
rect 3712 7584 3776 7588
rect 3792 7644 3856 7648
rect 3792 7588 3796 7644
rect 3796 7588 3852 7644
rect 3852 7588 3856 7644
rect 3792 7584 3856 7588
rect 3872 7644 3936 7648
rect 3872 7588 3876 7644
rect 3876 7588 3932 7644
rect 3932 7588 3936 7644
rect 3872 7584 3936 7588
rect 3952 7644 4016 7648
rect 3952 7588 3956 7644
rect 3956 7588 4012 7644
rect 4012 7588 4016 7644
rect 3952 7584 4016 7588
rect 5920 7644 5984 7648
rect 5920 7588 5924 7644
rect 5924 7588 5980 7644
rect 5980 7588 5984 7644
rect 5920 7584 5984 7588
rect 6000 7644 6064 7648
rect 6000 7588 6004 7644
rect 6004 7588 6060 7644
rect 6060 7588 6064 7644
rect 6000 7584 6064 7588
rect 6080 7644 6144 7648
rect 6080 7588 6084 7644
rect 6084 7588 6140 7644
rect 6140 7588 6144 7644
rect 6080 7584 6144 7588
rect 6160 7644 6224 7648
rect 6160 7588 6164 7644
rect 6164 7588 6220 7644
rect 6220 7588 6224 7644
rect 6160 7584 6224 7588
rect 8128 7644 8192 7648
rect 8128 7588 8132 7644
rect 8132 7588 8188 7644
rect 8188 7588 8192 7644
rect 8128 7584 8192 7588
rect 8208 7644 8272 7648
rect 8208 7588 8212 7644
rect 8212 7588 8268 7644
rect 8268 7588 8272 7644
rect 8208 7584 8272 7588
rect 8288 7644 8352 7648
rect 8288 7588 8292 7644
rect 8292 7588 8348 7644
rect 8348 7588 8352 7644
rect 8288 7584 8352 7588
rect 8368 7644 8432 7648
rect 8368 7588 8372 7644
rect 8372 7588 8428 7644
rect 8428 7588 8432 7644
rect 8368 7584 8432 7588
rect 2608 7100 2672 7104
rect 2608 7044 2612 7100
rect 2612 7044 2668 7100
rect 2668 7044 2672 7100
rect 2608 7040 2672 7044
rect 2688 7100 2752 7104
rect 2688 7044 2692 7100
rect 2692 7044 2748 7100
rect 2748 7044 2752 7100
rect 2688 7040 2752 7044
rect 2768 7100 2832 7104
rect 2768 7044 2772 7100
rect 2772 7044 2828 7100
rect 2828 7044 2832 7100
rect 2768 7040 2832 7044
rect 2848 7100 2912 7104
rect 2848 7044 2852 7100
rect 2852 7044 2908 7100
rect 2908 7044 2912 7100
rect 2848 7040 2912 7044
rect 4816 7100 4880 7104
rect 4816 7044 4820 7100
rect 4820 7044 4876 7100
rect 4876 7044 4880 7100
rect 4816 7040 4880 7044
rect 4896 7100 4960 7104
rect 4896 7044 4900 7100
rect 4900 7044 4956 7100
rect 4956 7044 4960 7100
rect 4896 7040 4960 7044
rect 4976 7100 5040 7104
rect 4976 7044 4980 7100
rect 4980 7044 5036 7100
rect 5036 7044 5040 7100
rect 4976 7040 5040 7044
rect 5056 7100 5120 7104
rect 5056 7044 5060 7100
rect 5060 7044 5116 7100
rect 5116 7044 5120 7100
rect 5056 7040 5120 7044
rect 7024 7100 7088 7104
rect 7024 7044 7028 7100
rect 7028 7044 7084 7100
rect 7084 7044 7088 7100
rect 7024 7040 7088 7044
rect 7104 7100 7168 7104
rect 7104 7044 7108 7100
rect 7108 7044 7164 7100
rect 7164 7044 7168 7100
rect 7104 7040 7168 7044
rect 7184 7100 7248 7104
rect 7184 7044 7188 7100
rect 7188 7044 7244 7100
rect 7244 7044 7248 7100
rect 7184 7040 7248 7044
rect 7264 7100 7328 7104
rect 7264 7044 7268 7100
rect 7268 7044 7324 7100
rect 7324 7044 7328 7100
rect 7264 7040 7328 7044
rect 9232 7100 9296 7104
rect 9232 7044 9236 7100
rect 9236 7044 9292 7100
rect 9292 7044 9296 7100
rect 9232 7040 9296 7044
rect 9312 7100 9376 7104
rect 9312 7044 9316 7100
rect 9316 7044 9372 7100
rect 9372 7044 9376 7100
rect 9312 7040 9376 7044
rect 9392 7100 9456 7104
rect 9392 7044 9396 7100
rect 9396 7044 9452 7100
rect 9452 7044 9456 7100
rect 9392 7040 9456 7044
rect 9472 7100 9536 7104
rect 9472 7044 9476 7100
rect 9476 7044 9532 7100
rect 9532 7044 9536 7100
rect 9472 7040 9536 7044
rect 1504 6556 1568 6560
rect 1504 6500 1508 6556
rect 1508 6500 1564 6556
rect 1564 6500 1568 6556
rect 1504 6496 1568 6500
rect 1584 6556 1648 6560
rect 1584 6500 1588 6556
rect 1588 6500 1644 6556
rect 1644 6500 1648 6556
rect 1584 6496 1648 6500
rect 1664 6556 1728 6560
rect 1664 6500 1668 6556
rect 1668 6500 1724 6556
rect 1724 6500 1728 6556
rect 1664 6496 1728 6500
rect 1744 6556 1808 6560
rect 1744 6500 1748 6556
rect 1748 6500 1804 6556
rect 1804 6500 1808 6556
rect 1744 6496 1808 6500
rect 3712 6556 3776 6560
rect 3712 6500 3716 6556
rect 3716 6500 3772 6556
rect 3772 6500 3776 6556
rect 3712 6496 3776 6500
rect 3792 6556 3856 6560
rect 3792 6500 3796 6556
rect 3796 6500 3852 6556
rect 3852 6500 3856 6556
rect 3792 6496 3856 6500
rect 3872 6556 3936 6560
rect 3872 6500 3876 6556
rect 3876 6500 3932 6556
rect 3932 6500 3936 6556
rect 3872 6496 3936 6500
rect 3952 6556 4016 6560
rect 3952 6500 3956 6556
rect 3956 6500 4012 6556
rect 4012 6500 4016 6556
rect 3952 6496 4016 6500
rect 5920 6556 5984 6560
rect 5920 6500 5924 6556
rect 5924 6500 5980 6556
rect 5980 6500 5984 6556
rect 5920 6496 5984 6500
rect 6000 6556 6064 6560
rect 6000 6500 6004 6556
rect 6004 6500 6060 6556
rect 6060 6500 6064 6556
rect 6000 6496 6064 6500
rect 6080 6556 6144 6560
rect 6080 6500 6084 6556
rect 6084 6500 6140 6556
rect 6140 6500 6144 6556
rect 6080 6496 6144 6500
rect 6160 6556 6224 6560
rect 6160 6500 6164 6556
rect 6164 6500 6220 6556
rect 6220 6500 6224 6556
rect 6160 6496 6224 6500
rect 8128 6556 8192 6560
rect 8128 6500 8132 6556
rect 8132 6500 8188 6556
rect 8188 6500 8192 6556
rect 8128 6496 8192 6500
rect 8208 6556 8272 6560
rect 8208 6500 8212 6556
rect 8212 6500 8268 6556
rect 8268 6500 8272 6556
rect 8208 6496 8272 6500
rect 8288 6556 8352 6560
rect 8288 6500 8292 6556
rect 8292 6500 8348 6556
rect 8348 6500 8352 6556
rect 8288 6496 8352 6500
rect 8368 6556 8432 6560
rect 8368 6500 8372 6556
rect 8372 6500 8428 6556
rect 8428 6500 8432 6556
rect 8368 6496 8432 6500
rect 2608 6012 2672 6016
rect 2608 5956 2612 6012
rect 2612 5956 2668 6012
rect 2668 5956 2672 6012
rect 2608 5952 2672 5956
rect 2688 6012 2752 6016
rect 2688 5956 2692 6012
rect 2692 5956 2748 6012
rect 2748 5956 2752 6012
rect 2688 5952 2752 5956
rect 2768 6012 2832 6016
rect 2768 5956 2772 6012
rect 2772 5956 2828 6012
rect 2828 5956 2832 6012
rect 2768 5952 2832 5956
rect 2848 6012 2912 6016
rect 2848 5956 2852 6012
rect 2852 5956 2908 6012
rect 2908 5956 2912 6012
rect 2848 5952 2912 5956
rect 4816 6012 4880 6016
rect 4816 5956 4820 6012
rect 4820 5956 4876 6012
rect 4876 5956 4880 6012
rect 4816 5952 4880 5956
rect 4896 6012 4960 6016
rect 4896 5956 4900 6012
rect 4900 5956 4956 6012
rect 4956 5956 4960 6012
rect 4896 5952 4960 5956
rect 4976 6012 5040 6016
rect 4976 5956 4980 6012
rect 4980 5956 5036 6012
rect 5036 5956 5040 6012
rect 4976 5952 5040 5956
rect 5056 6012 5120 6016
rect 5056 5956 5060 6012
rect 5060 5956 5116 6012
rect 5116 5956 5120 6012
rect 5056 5952 5120 5956
rect 7024 6012 7088 6016
rect 7024 5956 7028 6012
rect 7028 5956 7084 6012
rect 7084 5956 7088 6012
rect 7024 5952 7088 5956
rect 7104 6012 7168 6016
rect 7104 5956 7108 6012
rect 7108 5956 7164 6012
rect 7164 5956 7168 6012
rect 7104 5952 7168 5956
rect 7184 6012 7248 6016
rect 7184 5956 7188 6012
rect 7188 5956 7244 6012
rect 7244 5956 7248 6012
rect 7184 5952 7248 5956
rect 7264 6012 7328 6016
rect 7264 5956 7268 6012
rect 7268 5956 7324 6012
rect 7324 5956 7328 6012
rect 7264 5952 7328 5956
rect 9232 6012 9296 6016
rect 9232 5956 9236 6012
rect 9236 5956 9292 6012
rect 9292 5956 9296 6012
rect 9232 5952 9296 5956
rect 9312 6012 9376 6016
rect 9312 5956 9316 6012
rect 9316 5956 9372 6012
rect 9372 5956 9376 6012
rect 9312 5952 9376 5956
rect 9392 6012 9456 6016
rect 9392 5956 9396 6012
rect 9396 5956 9452 6012
rect 9452 5956 9456 6012
rect 9392 5952 9456 5956
rect 9472 6012 9536 6016
rect 9472 5956 9476 6012
rect 9476 5956 9532 6012
rect 9532 5956 9536 6012
rect 9472 5952 9536 5956
rect 1504 5468 1568 5472
rect 1504 5412 1508 5468
rect 1508 5412 1564 5468
rect 1564 5412 1568 5468
rect 1504 5408 1568 5412
rect 1584 5468 1648 5472
rect 1584 5412 1588 5468
rect 1588 5412 1644 5468
rect 1644 5412 1648 5468
rect 1584 5408 1648 5412
rect 1664 5468 1728 5472
rect 1664 5412 1668 5468
rect 1668 5412 1724 5468
rect 1724 5412 1728 5468
rect 1664 5408 1728 5412
rect 1744 5468 1808 5472
rect 1744 5412 1748 5468
rect 1748 5412 1804 5468
rect 1804 5412 1808 5468
rect 1744 5408 1808 5412
rect 3712 5468 3776 5472
rect 3712 5412 3716 5468
rect 3716 5412 3772 5468
rect 3772 5412 3776 5468
rect 3712 5408 3776 5412
rect 3792 5468 3856 5472
rect 3792 5412 3796 5468
rect 3796 5412 3852 5468
rect 3852 5412 3856 5468
rect 3792 5408 3856 5412
rect 3872 5468 3936 5472
rect 3872 5412 3876 5468
rect 3876 5412 3932 5468
rect 3932 5412 3936 5468
rect 3872 5408 3936 5412
rect 3952 5468 4016 5472
rect 3952 5412 3956 5468
rect 3956 5412 4012 5468
rect 4012 5412 4016 5468
rect 3952 5408 4016 5412
rect 5920 5468 5984 5472
rect 5920 5412 5924 5468
rect 5924 5412 5980 5468
rect 5980 5412 5984 5468
rect 5920 5408 5984 5412
rect 6000 5468 6064 5472
rect 6000 5412 6004 5468
rect 6004 5412 6060 5468
rect 6060 5412 6064 5468
rect 6000 5408 6064 5412
rect 6080 5468 6144 5472
rect 6080 5412 6084 5468
rect 6084 5412 6140 5468
rect 6140 5412 6144 5468
rect 6080 5408 6144 5412
rect 6160 5468 6224 5472
rect 6160 5412 6164 5468
rect 6164 5412 6220 5468
rect 6220 5412 6224 5468
rect 6160 5408 6224 5412
rect 8128 5468 8192 5472
rect 8128 5412 8132 5468
rect 8132 5412 8188 5468
rect 8188 5412 8192 5468
rect 8128 5408 8192 5412
rect 8208 5468 8272 5472
rect 8208 5412 8212 5468
rect 8212 5412 8268 5468
rect 8268 5412 8272 5468
rect 8208 5408 8272 5412
rect 8288 5468 8352 5472
rect 8288 5412 8292 5468
rect 8292 5412 8348 5468
rect 8348 5412 8352 5468
rect 8288 5408 8352 5412
rect 8368 5468 8432 5472
rect 8368 5412 8372 5468
rect 8372 5412 8428 5468
rect 8428 5412 8432 5468
rect 8368 5408 8432 5412
rect 2608 4924 2672 4928
rect 2608 4868 2612 4924
rect 2612 4868 2668 4924
rect 2668 4868 2672 4924
rect 2608 4864 2672 4868
rect 2688 4924 2752 4928
rect 2688 4868 2692 4924
rect 2692 4868 2748 4924
rect 2748 4868 2752 4924
rect 2688 4864 2752 4868
rect 2768 4924 2832 4928
rect 2768 4868 2772 4924
rect 2772 4868 2828 4924
rect 2828 4868 2832 4924
rect 2768 4864 2832 4868
rect 2848 4924 2912 4928
rect 2848 4868 2852 4924
rect 2852 4868 2908 4924
rect 2908 4868 2912 4924
rect 2848 4864 2912 4868
rect 4816 4924 4880 4928
rect 4816 4868 4820 4924
rect 4820 4868 4876 4924
rect 4876 4868 4880 4924
rect 4816 4864 4880 4868
rect 4896 4924 4960 4928
rect 4896 4868 4900 4924
rect 4900 4868 4956 4924
rect 4956 4868 4960 4924
rect 4896 4864 4960 4868
rect 4976 4924 5040 4928
rect 4976 4868 4980 4924
rect 4980 4868 5036 4924
rect 5036 4868 5040 4924
rect 4976 4864 5040 4868
rect 5056 4924 5120 4928
rect 5056 4868 5060 4924
rect 5060 4868 5116 4924
rect 5116 4868 5120 4924
rect 5056 4864 5120 4868
rect 7024 4924 7088 4928
rect 7024 4868 7028 4924
rect 7028 4868 7084 4924
rect 7084 4868 7088 4924
rect 7024 4864 7088 4868
rect 7104 4924 7168 4928
rect 7104 4868 7108 4924
rect 7108 4868 7164 4924
rect 7164 4868 7168 4924
rect 7104 4864 7168 4868
rect 7184 4924 7248 4928
rect 7184 4868 7188 4924
rect 7188 4868 7244 4924
rect 7244 4868 7248 4924
rect 7184 4864 7248 4868
rect 7264 4924 7328 4928
rect 7264 4868 7268 4924
rect 7268 4868 7324 4924
rect 7324 4868 7328 4924
rect 7264 4864 7328 4868
rect 9232 4924 9296 4928
rect 9232 4868 9236 4924
rect 9236 4868 9292 4924
rect 9292 4868 9296 4924
rect 9232 4864 9296 4868
rect 9312 4924 9376 4928
rect 9312 4868 9316 4924
rect 9316 4868 9372 4924
rect 9372 4868 9376 4924
rect 9312 4864 9376 4868
rect 9392 4924 9456 4928
rect 9392 4868 9396 4924
rect 9396 4868 9452 4924
rect 9452 4868 9456 4924
rect 9392 4864 9456 4868
rect 9472 4924 9536 4928
rect 9472 4868 9476 4924
rect 9476 4868 9532 4924
rect 9532 4868 9536 4924
rect 9472 4864 9536 4868
rect 1504 4380 1568 4384
rect 1504 4324 1508 4380
rect 1508 4324 1564 4380
rect 1564 4324 1568 4380
rect 1504 4320 1568 4324
rect 1584 4380 1648 4384
rect 1584 4324 1588 4380
rect 1588 4324 1644 4380
rect 1644 4324 1648 4380
rect 1584 4320 1648 4324
rect 1664 4380 1728 4384
rect 1664 4324 1668 4380
rect 1668 4324 1724 4380
rect 1724 4324 1728 4380
rect 1664 4320 1728 4324
rect 1744 4380 1808 4384
rect 1744 4324 1748 4380
rect 1748 4324 1804 4380
rect 1804 4324 1808 4380
rect 1744 4320 1808 4324
rect 3712 4380 3776 4384
rect 3712 4324 3716 4380
rect 3716 4324 3772 4380
rect 3772 4324 3776 4380
rect 3712 4320 3776 4324
rect 3792 4380 3856 4384
rect 3792 4324 3796 4380
rect 3796 4324 3852 4380
rect 3852 4324 3856 4380
rect 3792 4320 3856 4324
rect 3872 4380 3936 4384
rect 3872 4324 3876 4380
rect 3876 4324 3932 4380
rect 3932 4324 3936 4380
rect 3872 4320 3936 4324
rect 3952 4380 4016 4384
rect 3952 4324 3956 4380
rect 3956 4324 4012 4380
rect 4012 4324 4016 4380
rect 3952 4320 4016 4324
rect 5920 4380 5984 4384
rect 5920 4324 5924 4380
rect 5924 4324 5980 4380
rect 5980 4324 5984 4380
rect 5920 4320 5984 4324
rect 6000 4380 6064 4384
rect 6000 4324 6004 4380
rect 6004 4324 6060 4380
rect 6060 4324 6064 4380
rect 6000 4320 6064 4324
rect 6080 4380 6144 4384
rect 6080 4324 6084 4380
rect 6084 4324 6140 4380
rect 6140 4324 6144 4380
rect 6080 4320 6144 4324
rect 6160 4380 6224 4384
rect 6160 4324 6164 4380
rect 6164 4324 6220 4380
rect 6220 4324 6224 4380
rect 6160 4320 6224 4324
rect 8128 4380 8192 4384
rect 8128 4324 8132 4380
rect 8132 4324 8188 4380
rect 8188 4324 8192 4380
rect 8128 4320 8192 4324
rect 8208 4380 8272 4384
rect 8208 4324 8212 4380
rect 8212 4324 8268 4380
rect 8268 4324 8272 4380
rect 8208 4320 8272 4324
rect 8288 4380 8352 4384
rect 8288 4324 8292 4380
rect 8292 4324 8348 4380
rect 8348 4324 8352 4380
rect 8288 4320 8352 4324
rect 8368 4380 8432 4384
rect 8368 4324 8372 4380
rect 8372 4324 8428 4380
rect 8428 4324 8432 4380
rect 8368 4320 8432 4324
rect 2608 3836 2672 3840
rect 2608 3780 2612 3836
rect 2612 3780 2668 3836
rect 2668 3780 2672 3836
rect 2608 3776 2672 3780
rect 2688 3836 2752 3840
rect 2688 3780 2692 3836
rect 2692 3780 2748 3836
rect 2748 3780 2752 3836
rect 2688 3776 2752 3780
rect 2768 3836 2832 3840
rect 2768 3780 2772 3836
rect 2772 3780 2828 3836
rect 2828 3780 2832 3836
rect 2768 3776 2832 3780
rect 2848 3836 2912 3840
rect 2848 3780 2852 3836
rect 2852 3780 2908 3836
rect 2908 3780 2912 3836
rect 2848 3776 2912 3780
rect 4816 3836 4880 3840
rect 4816 3780 4820 3836
rect 4820 3780 4876 3836
rect 4876 3780 4880 3836
rect 4816 3776 4880 3780
rect 4896 3836 4960 3840
rect 4896 3780 4900 3836
rect 4900 3780 4956 3836
rect 4956 3780 4960 3836
rect 4896 3776 4960 3780
rect 4976 3836 5040 3840
rect 4976 3780 4980 3836
rect 4980 3780 5036 3836
rect 5036 3780 5040 3836
rect 4976 3776 5040 3780
rect 5056 3836 5120 3840
rect 5056 3780 5060 3836
rect 5060 3780 5116 3836
rect 5116 3780 5120 3836
rect 5056 3776 5120 3780
rect 7024 3836 7088 3840
rect 7024 3780 7028 3836
rect 7028 3780 7084 3836
rect 7084 3780 7088 3836
rect 7024 3776 7088 3780
rect 7104 3836 7168 3840
rect 7104 3780 7108 3836
rect 7108 3780 7164 3836
rect 7164 3780 7168 3836
rect 7104 3776 7168 3780
rect 7184 3836 7248 3840
rect 7184 3780 7188 3836
rect 7188 3780 7244 3836
rect 7244 3780 7248 3836
rect 7184 3776 7248 3780
rect 7264 3836 7328 3840
rect 7264 3780 7268 3836
rect 7268 3780 7324 3836
rect 7324 3780 7328 3836
rect 7264 3776 7328 3780
rect 9232 3836 9296 3840
rect 9232 3780 9236 3836
rect 9236 3780 9292 3836
rect 9292 3780 9296 3836
rect 9232 3776 9296 3780
rect 9312 3836 9376 3840
rect 9312 3780 9316 3836
rect 9316 3780 9372 3836
rect 9372 3780 9376 3836
rect 9312 3776 9376 3780
rect 9392 3836 9456 3840
rect 9392 3780 9396 3836
rect 9396 3780 9452 3836
rect 9452 3780 9456 3836
rect 9392 3776 9456 3780
rect 9472 3836 9536 3840
rect 9472 3780 9476 3836
rect 9476 3780 9532 3836
rect 9532 3780 9536 3836
rect 9472 3776 9536 3780
rect 1504 3292 1568 3296
rect 1504 3236 1508 3292
rect 1508 3236 1564 3292
rect 1564 3236 1568 3292
rect 1504 3232 1568 3236
rect 1584 3292 1648 3296
rect 1584 3236 1588 3292
rect 1588 3236 1644 3292
rect 1644 3236 1648 3292
rect 1584 3232 1648 3236
rect 1664 3292 1728 3296
rect 1664 3236 1668 3292
rect 1668 3236 1724 3292
rect 1724 3236 1728 3292
rect 1664 3232 1728 3236
rect 1744 3292 1808 3296
rect 1744 3236 1748 3292
rect 1748 3236 1804 3292
rect 1804 3236 1808 3292
rect 1744 3232 1808 3236
rect 3712 3292 3776 3296
rect 3712 3236 3716 3292
rect 3716 3236 3772 3292
rect 3772 3236 3776 3292
rect 3712 3232 3776 3236
rect 3792 3292 3856 3296
rect 3792 3236 3796 3292
rect 3796 3236 3852 3292
rect 3852 3236 3856 3292
rect 3792 3232 3856 3236
rect 3872 3292 3936 3296
rect 3872 3236 3876 3292
rect 3876 3236 3932 3292
rect 3932 3236 3936 3292
rect 3872 3232 3936 3236
rect 3952 3292 4016 3296
rect 3952 3236 3956 3292
rect 3956 3236 4012 3292
rect 4012 3236 4016 3292
rect 3952 3232 4016 3236
rect 5920 3292 5984 3296
rect 5920 3236 5924 3292
rect 5924 3236 5980 3292
rect 5980 3236 5984 3292
rect 5920 3232 5984 3236
rect 6000 3292 6064 3296
rect 6000 3236 6004 3292
rect 6004 3236 6060 3292
rect 6060 3236 6064 3292
rect 6000 3232 6064 3236
rect 6080 3292 6144 3296
rect 6080 3236 6084 3292
rect 6084 3236 6140 3292
rect 6140 3236 6144 3292
rect 6080 3232 6144 3236
rect 6160 3292 6224 3296
rect 6160 3236 6164 3292
rect 6164 3236 6220 3292
rect 6220 3236 6224 3292
rect 6160 3232 6224 3236
rect 8128 3292 8192 3296
rect 8128 3236 8132 3292
rect 8132 3236 8188 3292
rect 8188 3236 8192 3292
rect 8128 3232 8192 3236
rect 8208 3292 8272 3296
rect 8208 3236 8212 3292
rect 8212 3236 8268 3292
rect 8268 3236 8272 3292
rect 8208 3232 8272 3236
rect 8288 3292 8352 3296
rect 8288 3236 8292 3292
rect 8292 3236 8348 3292
rect 8348 3236 8352 3292
rect 8288 3232 8352 3236
rect 8368 3292 8432 3296
rect 8368 3236 8372 3292
rect 8372 3236 8428 3292
rect 8428 3236 8432 3292
rect 8368 3232 8432 3236
rect 2608 2748 2672 2752
rect 2608 2692 2612 2748
rect 2612 2692 2668 2748
rect 2668 2692 2672 2748
rect 2608 2688 2672 2692
rect 2688 2748 2752 2752
rect 2688 2692 2692 2748
rect 2692 2692 2748 2748
rect 2748 2692 2752 2748
rect 2688 2688 2752 2692
rect 2768 2748 2832 2752
rect 2768 2692 2772 2748
rect 2772 2692 2828 2748
rect 2828 2692 2832 2748
rect 2768 2688 2832 2692
rect 2848 2748 2912 2752
rect 2848 2692 2852 2748
rect 2852 2692 2908 2748
rect 2908 2692 2912 2748
rect 2848 2688 2912 2692
rect 4816 2748 4880 2752
rect 4816 2692 4820 2748
rect 4820 2692 4876 2748
rect 4876 2692 4880 2748
rect 4816 2688 4880 2692
rect 4896 2748 4960 2752
rect 4896 2692 4900 2748
rect 4900 2692 4956 2748
rect 4956 2692 4960 2748
rect 4896 2688 4960 2692
rect 4976 2748 5040 2752
rect 4976 2692 4980 2748
rect 4980 2692 5036 2748
rect 5036 2692 5040 2748
rect 4976 2688 5040 2692
rect 5056 2748 5120 2752
rect 5056 2692 5060 2748
rect 5060 2692 5116 2748
rect 5116 2692 5120 2748
rect 5056 2688 5120 2692
rect 7024 2748 7088 2752
rect 7024 2692 7028 2748
rect 7028 2692 7084 2748
rect 7084 2692 7088 2748
rect 7024 2688 7088 2692
rect 7104 2748 7168 2752
rect 7104 2692 7108 2748
rect 7108 2692 7164 2748
rect 7164 2692 7168 2748
rect 7104 2688 7168 2692
rect 7184 2748 7248 2752
rect 7184 2692 7188 2748
rect 7188 2692 7244 2748
rect 7244 2692 7248 2748
rect 7184 2688 7248 2692
rect 7264 2748 7328 2752
rect 7264 2692 7268 2748
rect 7268 2692 7324 2748
rect 7324 2692 7328 2748
rect 7264 2688 7328 2692
rect 9232 2748 9296 2752
rect 9232 2692 9236 2748
rect 9236 2692 9292 2748
rect 9292 2692 9296 2748
rect 9232 2688 9296 2692
rect 9312 2748 9376 2752
rect 9312 2692 9316 2748
rect 9316 2692 9372 2748
rect 9372 2692 9376 2748
rect 9312 2688 9376 2692
rect 9392 2748 9456 2752
rect 9392 2692 9396 2748
rect 9396 2692 9452 2748
rect 9452 2692 9456 2748
rect 9392 2688 9456 2692
rect 9472 2748 9536 2752
rect 9472 2692 9476 2748
rect 9476 2692 9532 2748
rect 9532 2692 9536 2748
rect 9472 2688 9536 2692
rect 1504 2204 1568 2208
rect 1504 2148 1508 2204
rect 1508 2148 1564 2204
rect 1564 2148 1568 2204
rect 1504 2144 1568 2148
rect 1584 2204 1648 2208
rect 1584 2148 1588 2204
rect 1588 2148 1644 2204
rect 1644 2148 1648 2204
rect 1584 2144 1648 2148
rect 1664 2204 1728 2208
rect 1664 2148 1668 2204
rect 1668 2148 1724 2204
rect 1724 2148 1728 2204
rect 1664 2144 1728 2148
rect 1744 2204 1808 2208
rect 1744 2148 1748 2204
rect 1748 2148 1804 2204
rect 1804 2148 1808 2204
rect 1744 2144 1808 2148
rect 3712 2204 3776 2208
rect 3712 2148 3716 2204
rect 3716 2148 3772 2204
rect 3772 2148 3776 2204
rect 3712 2144 3776 2148
rect 3792 2204 3856 2208
rect 3792 2148 3796 2204
rect 3796 2148 3852 2204
rect 3852 2148 3856 2204
rect 3792 2144 3856 2148
rect 3872 2204 3936 2208
rect 3872 2148 3876 2204
rect 3876 2148 3932 2204
rect 3932 2148 3936 2204
rect 3872 2144 3936 2148
rect 3952 2204 4016 2208
rect 3952 2148 3956 2204
rect 3956 2148 4012 2204
rect 4012 2148 4016 2204
rect 3952 2144 4016 2148
rect 5920 2204 5984 2208
rect 5920 2148 5924 2204
rect 5924 2148 5980 2204
rect 5980 2148 5984 2204
rect 5920 2144 5984 2148
rect 6000 2204 6064 2208
rect 6000 2148 6004 2204
rect 6004 2148 6060 2204
rect 6060 2148 6064 2204
rect 6000 2144 6064 2148
rect 6080 2204 6144 2208
rect 6080 2148 6084 2204
rect 6084 2148 6140 2204
rect 6140 2148 6144 2204
rect 6080 2144 6144 2148
rect 6160 2204 6224 2208
rect 6160 2148 6164 2204
rect 6164 2148 6220 2204
rect 6220 2148 6224 2204
rect 6160 2144 6224 2148
rect 8128 2204 8192 2208
rect 8128 2148 8132 2204
rect 8132 2148 8188 2204
rect 8188 2148 8192 2204
rect 8128 2144 8192 2148
rect 8208 2204 8272 2208
rect 8208 2148 8212 2204
rect 8212 2148 8268 2204
rect 8268 2148 8272 2204
rect 8208 2144 8272 2148
rect 8288 2204 8352 2208
rect 8288 2148 8292 2204
rect 8292 2148 8348 2204
rect 8348 2148 8352 2204
rect 8288 2144 8352 2148
rect 8368 2204 8432 2208
rect 8368 2148 8372 2204
rect 8372 2148 8428 2204
rect 8428 2148 8432 2204
rect 8368 2144 8432 2148
rect 2608 1660 2672 1664
rect 2608 1604 2612 1660
rect 2612 1604 2668 1660
rect 2668 1604 2672 1660
rect 2608 1600 2672 1604
rect 2688 1660 2752 1664
rect 2688 1604 2692 1660
rect 2692 1604 2748 1660
rect 2748 1604 2752 1660
rect 2688 1600 2752 1604
rect 2768 1660 2832 1664
rect 2768 1604 2772 1660
rect 2772 1604 2828 1660
rect 2828 1604 2832 1660
rect 2768 1600 2832 1604
rect 2848 1660 2912 1664
rect 2848 1604 2852 1660
rect 2852 1604 2908 1660
rect 2908 1604 2912 1660
rect 2848 1600 2912 1604
rect 4816 1660 4880 1664
rect 4816 1604 4820 1660
rect 4820 1604 4876 1660
rect 4876 1604 4880 1660
rect 4816 1600 4880 1604
rect 4896 1660 4960 1664
rect 4896 1604 4900 1660
rect 4900 1604 4956 1660
rect 4956 1604 4960 1660
rect 4896 1600 4960 1604
rect 4976 1660 5040 1664
rect 4976 1604 4980 1660
rect 4980 1604 5036 1660
rect 5036 1604 5040 1660
rect 4976 1600 5040 1604
rect 5056 1660 5120 1664
rect 5056 1604 5060 1660
rect 5060 1604 5116 1660
rect 5116 1604 5120 1660
rect 5056 1600 5120 1604
rect 7024 1660 7088 1664
rect 7024 1604 7028 1660
rect 7028 1604 7084 1660
rect 7084 1604 7088 1660
rect 7024 1600 7088 1604
rect 7104 1660 7168 1664
rect 7104 1604 7108 1660
rect 7108 1604 7164 1660
rect 7164 1604 7168 1660
rect 7104 1600 7168 1604
rect 7184 1660 7248 1664
rect 7184 1604 7188 1660
rect 7188 1604 7244 1660
rect 7244 1604 7248 1660
rect 7184 1600 7248 1604
rect 7264 1660 7328 1664
rect 7264 1604 7268 1660
rect 7268 1604 7324 1660
rect 7324 1604 7328 1660
rect 7264 1600 7328 1604
rect 9232 1660 9296 1664
rect 9232 1604 9236 1660
rect 9236 1604 9292 1660
rect 9292 1604 9296 1660
rect 9232 1600 9296 1604
rect 9312 1660 9376 1664
rect 9312 1604 9316 1660
rect 9316 1604 9372 1660
rect 9372 1604 9376 1660
rect 9312 1600 9376 1604
rect 9392 1660 9456 1664
rect 9392 1604 9396 1660
rect 9396 1604 9452 1660
rect 9452 1604 9456 1660
rect 9392 1600 9456 1604
rect 9472 1660 9536 1664
rect 9472 1604 9476 1660
rect 9476 1604 9532 1660
rect 9532 1604 9536 1660
rect 9472 1600 9536 1604
rect 1504 1116 1568 1120
rect 1504 1060 1508 1116
rect 1508 1060 1564 1116
rect 1564 1060 1568 1116
rect 1504 1056 1568 1060
rect 1584 1116 1648 1120
rect 1584 1060 1588 1116
rect 1588 1060 1644 1116
rect 1644 1060 1648 1116
rect 1584 1056 1648 1060
rect 1664 1116 1728 1120
rect 1664 1060 1668 1116
rect 1668 1060 1724 1116
rect 1724 1060 1728 1116
rect 1664 1056 1728 1060
rect 1744 1116 1808 1120
rect 1744 1060 1748 1116
rect 1748 1060 1804 1116
rect 1804 1060 1808 1116
rect 1744 1056 1808 1060
rect 3712 1116 3776 1120
rect 3712 1060 3716 1116
rect 3716 1060 3772 1116
rect 3772 1060 3776 1116
rect 3712 1056 3776 1060
rect 3792 1116 3856 1120
rect 3792 1060 3796 1116
rect 3796 1060 3852 1116
rect 3852 1060 3856 1116
rect 3792 1056 3856 1060
rect 3872 1116 3936 1120
rect 3872 1060 3876 1116
rect 3876 1060 3932 1116
rect 3932 1060 3936 1116
rect 3872 1056 3936 1060
rect 3952 1116 4016 1120
rect 3952 1060 3956 1116
rect 3956 1060 4012 1116
rect 4012 1060 4016 1116
rect 3952 1056 4016 1060
rect 5920 1116 5984 1120
rect 5920 1060 5924 1116
rect 5924 1060 5980 1116
rect 5980 1060 5984 1116
rect 5920 1056 5984 1060
rect 6000 1116 6064 1120
rect 6000 1060 6004 1116
rect 6004 1060 6060 1116
rect 6060 1060 6064 1116
rect 6000 1056 6064 1060
rect 6080 1116 6144 1120
rect 6080 1060 6084 1116
rect 6084 1060 6140 1116
rect 6140 1060 6144 1116
rect 6080 1056 6144 1060
rect 6160 1116 6224 1120
rect 6160 1060 6164 1116
rect 6164 1060 6220 1116
rect 6220 1060 6224 1116
rect 6160 1056 6224 1060
rect 8128 1116 8192 1120
rect 8128 1060 8132 1116
rect 8132 1060 8188 1116
rect 8188 1060 8192 1116
rect 8128 1056 8192 1060
rect 8208 1116 8272 1120
rect 8208 1060 8212 1116
rect 8212 1060 8268 1116
rect 8268 1060 8272 1116
rect 8208 1056 8272 1060
rect 8288 1116 8352 1120
rect 8288 1060 8292 1116
rect 8292 1060 8348 1116
rect 8348 1060 8352 1116
rect 8288 1056 8352 1060
rect 8368 1116 8432 1120
rect 8368 1060 8372 1116
rect 8372 1060 8428 1116
rect 8428 1060 8432 1116
rect 8368 1056 8432 1060
rect 2608 572 2672 576
rect 2608 516 2612 572
rect 2612 516 2668 572
rect 2668 516 2672 572
rect 2608 512 2672 516
rect 2688 572 2752 576
rect 2688 516 2692 572
rect 2692 516 2748 572
rect 2748 516 2752 572
rect 2688 512 2752 516
rect 2768 572 2832 576
rect 2768 516 2772 572
rect 2772 516 2828 572
rect 2828 516 2832 572
rect 2768 512 2832 516
rect 2848 572 2912 576
rect 2848 516 2852 572
rect 2852 516 2908 572
rect 2908 516 2912 572
rect 2848 512 2912 516
rect 4816 572 4880 576
rect 4816 516 4820 572
rect 4820 516 4876 572
rect 4876 516 4880 572
rect 4816 512 4880 516
rect 4896 572 4960 576
rect 4896 516 4900 572
rect 4900 516 4956 572
rect 4956 516 4960 572
rect 4896 512 4960 516
rect 4976 572 5040 576
rect 4976 516 4980 572
rect 4980 516 5036 572
rect 5036 516 5040 572
rect 4976 512 5040 516
rect 5056 572 5120 576
rect 5056 516 5060 572
rect 5060 516 5116 572
rect 5116 516 5120 572
rect 5056 512 5120 516
rect 7024 572 7088 576
rect 7024 516 7028 572
rect 7028 516 7084 572
rect 7084 516 7088 572
rect 7024 512 7088 516
rect 7104 572 7168 576
rect 7104 516 7108 572
rect 7108 516 7164 572
rect 7164 516 7168 572
rect 7104 512 7168 516
rect 7184 572 7248 576
rect 7184 516 7188 572
rect 7188 516 7244 572
rect 7244 516 7248 572
rect 7184 512 7248 516
rect 7264 572 7328 576
rect 7264 516 7268 572
rect 7268 516 7324 572
rect 7324 516 7328 572
rect 7264 512 7328 516
rect 9232 572 9296 576
rect 9232 516 9236 572
rect 9236 516 9292 572
rect 9292 516 9296 572
rect 9232 512 9296 516
rect 9312 572 9376 576
rect 9312 516 9316 572
rect 9316 516 9372 572
rect 9372 516 9376 572
rect 9312 512 9376 516
rect 9392 572 9456 576
rect 9392 516 9396 572
rect 9396 516 9452 572
rect 9452 516 9456 572
rect 9392 512 9456 516
rect 9472 572 9536 576
rect 9472 516 9476 572
rect 9476 516 9532 572
rect 9532 516 9536 572
rect 9472 512 9536 516
<< metal4 >>
rect 1496 8736 1816 9296
rect 1496 8672 1504 8736
rect 1568 8672 1584 8736
rect 1648 8672 1664 8736
rect 1728 8672 1744 8736
rect 1808 8672 1816 8736
rect 1496 7648 1816 8672
rect 1496 7584 1504 7648
rect 1568 7584 1584 7648
rect 1648 7584 1664 7648
rect 1728 7584 1744 7648
rect 1808 7584 1816 7648
rect 1496 6560 1816 7584
rect 1496 6496 1504 6560
rect 1568 6496 1584 6560
rect 1648 6496 1664 6560
rect 1728 6496 1744 6560
rect 1808 6496 1816 6560
rect 1496 5472 1816 6496
rect 1496 5408 1504 5472
rect 1568 5408 1584 5472
rect 1648 5408 1664 5472
rect 1728 5408 1744 5472
rect 1808 5408 1816 5472
rect 1496 4384 1816 5408
rect 1496 4320 1504 4384
rect 1568 4320 1584 4384
rect 1648 4320 1664 4384
rect 1728 4320 1744 4384
rect 1808 4320 1816 4384
rect 1496 3296 1816 4320
rect 1496 3232 1504 3296
rect 1568 3232 1584 3296
rect 1648 3232 1664 3296
rect 1728 3232 1744 3296
rect 1808 3232 1816 3296
rect 1496 2208 1816 3232
rect 1496 2144 1504 2208
rect 1568 2144 1584 2208
rect 1648 2144 1664 2208
rect 1728 2144 1744 2208
rect 1808 2144 1816 2208
rect 1496 1120 1816 2144
rect 1496 1056 1504 1120
rect 1568 1056 1584 1120
rect 1648 1056 1664 1120
rect 1728 1056 1744 1120
rect 1808 1056 1816 1120
rect 1496 496 1816 1056
rect 2600 9280 2920 9296
rect 2600 9216 2608 9280
rect 2672 9216 2688 9280
rect 2752 9216 2768 9280
rect 2832 9216 2848 9280
rect 2912 9216 2920 9280
rect 2600 8192 2920 9216
rect 2600 8128 2608 8192
rect 2672 8128 2688 8192
rect 2752 8128 2768 8192
rect 2832 8128 2848 8192
rect 2912 8128 2920 8192
rect 2600 7104 2920 8128
rect 2600 7040 2608 7104
rect 2672 7040 2688 7104
rect 2752 7040 2768 7104
rect 2832 7040 2848 7104
rect 2912 7040 2920 7104
rect 2600 6016 2920 7040
rect 2600 5952 2608 6016
rect 2672 5952 2688 6016
rect 2752 5952 2768 6016
rect 2832 5952 2848 6016
rect 2912 5952 2920 6016
rect 2600 4928 2920 5952
rect 2600 4864 2608 4928
rect 2672 4864 2688 4928
rect 2752 4864 2768 4928
rect 2832 4864 2848 4928
rect 2912 4864 2920 4928
rect 2600 3840 2920 4864
rect 2600 3776 2608 3840
rect 2672 3776 2688 3840
rect 2752 3776 2768 3840
rect 2832 3776 2848 3840
rect 2912 3776 2920 3840
rect 2600 2752 2920 3776
rect 2600 2688 2608 2752
rect 2672 2688 2688 2752
rect 2752 2688 2768 2752
rect 2832 2688 2848 2752
rect 2912 2688 2920 2752
rect 2600 1664 2920 2688
rect 2600 1600 2608 1664
rect 2672 1600 2688 1664
rect 2752 1600 2768 1664
rect 2832 1600 2848 1664
rect 2912 1600 2920 1664
rect 2600 576 2920 1600
rect 2600 512 2608 576
rect 2672 512 2688 576
rect 2752 512 2768 576
rect 2832 512 2848 576
rect 2912 512 2920 576
rect 2600 496 2920 512
rect 3704 8736 4024 9296
rect 3704 8672 3712 8736
rect 3776 8672 3792 8736
rect 3856 8672 3872 8736
rect 3936 8672 3952 8736
rect 4016 8672 4024 8736
rect 3704 7648 4024 8672
rect 3704 7584 3712 7648
rect 3776 7584 3792 7648
rect 3856 7584 3872 7648
rect 3936 7584 3952 7648
rect 4016 7584 4024 7648
rect 3704 6560 4024 7584
rect 3704 6496 3712 6560
rect 3776 6496 3792 6560
rect 3856 6496 3872 6560
rect 3936 6496 3952 6560
rect 4016 6496 4024 6560
rect 3704 5472 4024 6496
rect 3704 5408 3712 5472
rect 3776 5408 3792 5472
rect 3856 5408 3872 5472
rect 3936 5408 3952 5472
rect 4016 5408 4024 5472
rect 3704 4384 4024 5408
rect 3704 4320 3712 4384
rect 3776 4320 3792 4384
rect 3856 4320 3872 4384
rect 3936 4320 3952 4384
rect 4016 4320 4024 4384
rect 3704 3296 4024 4320
rect 3704 3232 3712 3296
rect 3776 3232 3792 3296
rect 3856 3232 3872 3296
rect 3936 3232 3952 3296
rect 4016 3232 4024 3296
rect 3704 2208 4024 3232
rect 3704 2144 3712 2208
rect 3776 2144 3792 2208
rect 3856 2144 3872 2208
rect 3936 2144 3952 2208
rect 4016 2144 4024 2208
rect 3704 1120 4024 2144
rect 3704 1056 3712 1120
rect 3776 1056 3792 1120
rect 3856 1056 3872 1120
rect 3936 1056 3952 1120
rect 4016 1056 4024 1120
rect 3704 496 4024 1056
rect 4808 9280 5128 9296
rect 4808 9216 4816 9280
rect 4880 9216 4896 9280
rect 4960 9216 4976 9280
rect 5040 9216 5056 9280
rect 5120 9216 5128 9280
rect 4808 8192 5128 9216
rect 4808 8128 4816 8192
rect 4880 8128 4896 8192
rect 4960 8128 4976 8192
rect 5040 8128 5056 8192
rect 5120 8128 5128 8192
rect 4808 7104 5128 8128
rect 4808 7040 4816 7104
rect 4880 7040 4896 7104
rect 4960 7040 4976 7104
rect 5040 7040 5056 7104
rect 5120 7040 5128 7104
rect 4808 6016 5128 7040
rect 4808 5952 4816 6016
rect 4880 5952 4896 6016
rect 4960 5952 4976 6016
rect 5040 5952 5056 6016
rect 5120 5952 5128 6016
rect 4808 4928 5128 5952
rect 4808 4864 4816 4928
rect 4880 4864 4896 4928
rect 4960 4864 4976 4928
rect 5040 4864 5056 4928
rect 5120 4864 5128 4928
rect 4808 3840 5128 4864
rect 4808 3776 4816 3840
rect 4880 3776 4896 3840
rect 4960 3776 4976 3840
rect 5040 3776 5056 3840
rect 5120 3776 5128 3840
rect 4808 2752 5128 3776
rect 4808 2688 4816 2752
rect 4880 2688 4896 2752
rect 4960 2688 4976 2752
rect 5040 2688 5056 2752
rect 5120 2688 5128 2752
rect 4808 1664 5128 2688
rect 4808 1600 4816 1664
rect 4880 1600 4896 1664
rect 4960 1600 4976 1664
rect 5040 1600 5056 1664
rect 5120 1600 5128 1664
rect 4808 576 5128 1600
rect 4808 512 4816 576
rect 4880 512 4896 576
rect 4960 512 4976 576
rect 5040 512 5056 576
rect 5120 512 5128 576
rect 4808 496 5128 512
rect 5912 8736 6232 9296
rect 5912 8672 5920 8736
rect 5984 8672 6000 8736
rect 6064 8672 6080 8736
rect 6144 8672 6160 8736
rect 6224 8672 6232 8736
rect 5912 7648 6232 8672
rect 5912 7584 5920 7648
rect 5984 7584 6000 7648
rect 6064 7584 6080 7648
rect 6144 7584 6160 7648
rect 6224 7584 6232 7648
rect 5912 6560 6232 7584
rect 5912 6496 5920 6560
rect 5984 6496 6000 6560
rect 6064 6496 6080 6560
rect 6144 6496 6160 6560
rect 6224 6496 6232 6560
rect 5912 5472 6232 6496
rect 5912 5408 5920 5472
rect 5984 5408 6000 5472
rect 6064 5408 6080 5472
rect 6144 5408 6160 5472
rect 6224 5408 6232 5472
rect 5912 4384 6232 5408
rect 5912 4320 5920 4384
rect 5984 4320 6000 4384
rect 6064 4320 6080 4384
rect 6144 4320 6160 4384
rect 6224 4320 6232 4384
rect 5912 3296 6232 4320
rect 5912 3232 5920 3296
rect 5984 3232 6000 3296
rect 6064 3232 6080 3296
rect 6144 3232 6160 3296
rect 6224 3232 6232 3296
rect 5912 2208 6232 3232
rect 5912 2144 5920 2208
rect 5984 2144 6000 2208
rect 6064 2144 6080 2208
rect 6144 2144 6160 2208
rect 6224 2144 6232 2208
rect 5912 1120 6232 2144
rect 5912 1056 5920 1120
rect 5984 1056 6000 1120
rect 6064 1056 6080 1120
rect 6144 1056 6160 1120
rect 6224 1056 6232 1120
rect 5912 496 6232 1056
rect 7016 9280 7336 9296
rect 7016 9216 7024 9280
rect 7088 9216 7104 9280
rect 7168 9216 7184 9280
rect 7248 9216 7264 9280
rect 7328 9216 7336 9280
rect 7016 8192 7336 9216
rect 7016 8128 7024 8192
rect 7088 8128 7104 8192
rect 7168 8128 7184 8192
rect 7248 8128 7264 8192
rect 7328 8128 7336 8192
rect 7016 7104 7336 8128
rect 7016 7040 7024 7104
rect 7088 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7336 7104
rect 7016 6016 7336 7040
rect 7016 5952 7024 6016
rect 7088 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7336 6016
rect 7016 4928 7336 5952
rect 7016 4864 7024 4928
rect 7088 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7336 4928
rect 7016 3840 7336 4864
rect 7016 3776 7024 3840
rect 7088 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7336 3840
rect 7016 2752 7336 3776
rect 7016 2688 7024 2752
rect 7088 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7336 2752
rect 7016 1664 7336 2688
rect 7016 1600 7024 1664
rect 7088 1600 7104 1664
rect 7168 1600 7184 1664
rect 7248 1600 7264 1664
rect 7328 1600 7336 1664
rect 7016 576 7336 1600
rect 7016 512 7024 576
rect 7088 512 7104 576
rect 7168 512 7184 576
rect 7248 512 7264 576
rect 7328 512 7336 576
rect 7016 496 7336 512
rect 8120 8736 8440 9296
rect 8120 8672 8128 8736
rect 8192 8672 8208 8736
rect 8272 8672 8288 8736
rect 8352 8672 8368 8736
rect 8432 8672 8440 8736
rect 8120 7648 8440 8672
rect 8120 7584 8128 7648
rect 8192 7584 8208 7648
rect 8272 7584 8288 7648
rect 8352 7584 8368 7648
rect 8432 7584 8440 7648
rect 8120 6560 8440 7584
rect 8120 6496 8128 6560
rect 8192 6496 8208 6560
rect 8272 6496 8288 6560
rect 8352 6496 8368 6560
rect 8432 6496 8440 6560
rect 8120 5472 8440 6496
rect 8120 5408 8128 5472
rect 8192 5408 8208 5472
rect 8272 5408 8288 5472
rect 8352 5408 8368 5472
rect 8432 5408 8440 5472
rect 8120 4384 8440 5408
rect 8120 4320 8128 4384
rect 8192 4320 8208 4384
rect 8272 4320 8288 4384
rect 8352 4320 8368 4384
rect 8432 4320 8440 4384
rect 8120 3296 8440 4320
rect 8120 3232 8128 3296
rect 8192 3232 8208 3296
rect 8272 3232 8288 3296
rect 8352 3232 8368 3296
rect 8432 3232 8440 3296
rect 8120 2208 8440 3232
rect 8120 2144 8128 2208
rect 8192 2144 8208 2208
rect 8272 2144 8288 2208
rect 8352 2144 8368 2208
rect 8432 2144 8440 2208
rect 8120 1120 8440 2144
rect 8120 1056 8128 1120
rect 8192 1056 8208 1120
rect 8272 1056 8288 1120
rect 8352 1056 8368 1120
rect 8432 1056 8440 1120
rect 8120 496 8440 1056
rect 9224 9280 9544 9296
rect 9224 9216 9232 9280
rect 9296 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9544 9280
rect 9224 8192 9544 9216
rect 9224 8128 9232 8192
rect 9296 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9544 8192
rect 9224 7104 9544 8128
rect 9224 7040 9232 7104
rect 9296 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9544 7104
rect 9224 6016 9544 7040
rect 9224 5952 9232 6016
rect 9296 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9544 6016
rect 9224 4928 9544 5952
rect 9224 4864 9232 4928
rect 9296 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9544 4928
rect 9224 3840 9544 4864
rect 9224 3776 9232 3840
rect 9296 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9544 3840
rect 9224 2752 9544 3776
rect 9224 2688 9232 2752
rect 9296 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9544 2752
rect 9224 1664 9544 2688
rect 9224 1600 9232 1664
rect 9296 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9544 1664
rect 9224 576 9544 1600
rect 9224 512 9232 576
rect 9296 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9544 576
rect 9224 496 9544 512
use sky130_fd_sc_hd__inv_2  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8832 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6808 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2760 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2576 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _16_
timestamp 1704896540
transform -1 0 3128 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 1704896540
transform -1 0 4232 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6532 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _20_
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23__2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6992 0 -1 1632
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_4  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8004 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _25_
timestamp 1704896540
transform -1 0 4324 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _26_
timestamp 1704896540
transform 1 0 3496 0 1 544
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _27_
timestamp 1704896540
transform 1 0 4876 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6716 0 1 1632
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 4508 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 6440 0 1 544
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2300 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1704896540
transform 1 0 8740 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_68
timestamp 1704896540
transform 1 0 6808 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_19
timestamp 1704896540
transform 1 0 2300 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_46
timestamp 1704896540
transform 1 0 4784 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_67
timestamp 1704896540
transform 1 0 6716 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_73
timestamp 1704896540
transform 1 0 7268 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_43
timestamp 1704896540
transform 1 0 4508 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_61
timestamp 1704896540
transform 1 0 6164 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_89
timestamp 1704896540
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_66
timestamp 1704896540
transform 1 0 6624 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_78
timestamp 1704896540
transform 1 0 7728 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_29
timestamp 1704896540
transform 1 0 3220 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_41
timestamp 1704896540
transform 1 0 4324 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1704896540
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_85
timestamp 1704896540
transform 1 0 8372 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9108 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 8740 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform -1 0 5060 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 3956 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 2392 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform 1 0 8832 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_16
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 9384 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_17
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 9384 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_18
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 9384 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_19
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_20
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 9384 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_21
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 9384 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_22
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 9384 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_23
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 9384 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_24
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 9384 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_25
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 9384 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_26
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 9384 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_27
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 9384 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_28
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 9384 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_29
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 9384 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_30
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_31
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 9384 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_35
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_38
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_39
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_40
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_41
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_42
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_43
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_44
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_45
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_46
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_47
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_48
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_49
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_50
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_51
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_52
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_53
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_54
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_55
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_56
timestamp 1704896540
transform 1 0 3128 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_57
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1704896540
transform 1 0 8280 0 -1 9248
box -38 -48 130 592
<< labels >>
rlabel metal2 s 5048 9248 5048 9248 4 VGND
rlabel metal1 s 4968 8704 4968 8704 4 VPWR
rlabel metal1 s 8747 1462 8747 1462 4 _00_
rlabel metal2 s 8602 1870 8602 1870 4 _01_
rlabel metal2 s 2530 1700 2530 1700 4 _02_
rlabel metal1 s 4048 782 4048 782 4 _03_
rlabel metal1 s 5244 986 5244 986 4 _04_
rlabel metal2 s 2346 1190 2346 1190 4 _05_
rlabel metal1 s 4002 1836 4002 1836 4 _06_
rlabel metal1 s 4922 1530 4922 1530 4 _07_
rlabel metal1 s 5934 1190 5934 1190 4 _08_
rlabel metal1 s 5658 986 5658 986 4 _09_
rlabel metal1 s 5520 782 5520 782 4 _10_
rlabel metal2 s 7498 1078 7498 1078 4 clk
rlabel metal1 s 5934 1734 5934 1734 4 clknet_0_clk
rlabel metal1 s 3680 2618 3680 2618 4 clknet_1_0__leaf_clk
rlabel metal2 s 7958 1700 7958 1700 4 clknet_1_1__leaf_clk
rlabel metal1 s 1702 646 1702 646 4 count[0]
rlabel metal1 s 2484 782 2484 782 4 count[1]
rlabel metal1 s 4738 646 4738 646 4 count[2]
rlabel metal2 s 5842 2074 5842 2074 4 count[3]
rlabel metal2 s 9154 568 9154 568 4 n_rst
rlabel metal2 s 8878 1190 8878 1190 4 net1
rlabel metal1 s 7360 1462 7360 1462 4 net2
rlabel metal2 s 6762 1156 6762 1156 4 net3
rlabel metal1 s 7866 2482 7866 2482 4 net4
rlabel metal1 s 3082 680 3082 680 4 net5
rlabel metal1 s 2162 1428 2162 1428 4 net6
rlabel metal1 s 3542 1394 3542 1394 4 net7
rlabel metal1 s 6302 1292 6302 1292 4 rst
flabel metal4 s 9224 496 9544 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7016 496 7336 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4808 496 5128 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2600 496 2920 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8120 496 8440 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5912 496 6232 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3704 496 4024 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1496 496 1816 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 7470 0 7526 400 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 846 0 902 400 0 FreeSans 280 90 0 0 count[0]
port 4 nsew
flabel metal2 s 2502 0 2558 400 0 FreeSans 280 90 0 0 count[1]
port 5 nsew
flabel metal2 s 4158 0 4214 400 0 FreeSans 280 90 0 0 count[2]
port 6 nsew
flabel metal2 s 5814 0 5870 400 0 FreeSans 280 90 0 0 count[3]
port 7 nsew
flabel metal2 s 9126 0 9182 400 0 FreeSans 280 90 0 0 n_rst
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string GDS_END 242986
string GDS_FILE ../gds/count_macro.gds
string GDS_START 113546
<< end >>
